// This is the unpowered netlist.
module serv_2 (io_in,
    io_oeb,
    io_out);
 input [4:0] io_in;
 output [4:0] io_oeb;
 output [4:0] io_out;

 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire _04725_;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire _04785_;
 wire _04786_;
 wire _04787_;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire _04809_;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire _04818_;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire \u_arbiter.i_wb_cpu_ack ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[10] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[11] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[12] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[13] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[14] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[15] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[16] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[17] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[18] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[19] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[20] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[21] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[22] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[23] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[24] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[25] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[26] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[27] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[28] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[29] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[2] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[30] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[31] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[3] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[4] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[5] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[6] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[7] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[8] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[9] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[0] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[10] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[11] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[12] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[13] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[14] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[15] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[16] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[17] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[18] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[19] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[1] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[20] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[21] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[22] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[23] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[24] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[25] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[26] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[27] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[28] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[29] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[2] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[30] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[31] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[3] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[4] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[5] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[6] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[7] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[8] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[9] ;
 wire \u_arbiter.i_wb_cpu_dbus_we ;
 wire \u_arbiter.i_wb_cpu_ibus_adr[0] ;
 wire \u_arbiter.i_wb_cpu_ibus_adr[1] ;
 wire \u_arbiter.i_wb_cpu_rdt[0] ;
 wire \u_arbiter.i_wb_cpu_rdt[10] ;
 wire \u_arbiter.i_wb_cpu_rdt[11] ;
 wire \u_arbiter.i_wb_cpu_rdt[12] ;
 wire \u_arbiter.i_wb_cpu_rdt[13] ;
 wire \u_arbiter.i_wb_cpu_rdt[14] ;
 wire \u_arbiter.i_wb_cpu_rdt[15] ;
 wire \u_arbiter.i_wb_cpu_rdt[16] ;
 wire \u_arbiter.i_wb_cpu_rdt[17] ;
 wire \u_arbiter.i_wb_cpu_rdt[18] ;
 wire \u_arbiter.i_wb_cpu_rdt[19] ;
 wire \u_arbiter.i_wb_cpu_rdt[1] ;
 wire \u_arbiter.i_wb_cpu_rdt[20] ;
 wire \u_arbiter.i_wb_cpu_rdt[21] ;
 wire \u_arbiter.i_wb_cpu_rdt[22] ;
 wire \u_arbiter.i_wb_cpu_rdt[23] ;
 wire \u_arbiter.i_wb_cpu_rdt[24] ;
 wire \u_arbiter.i_wb_cpu_rdt[25] ;
 wire \u_arbiter.i_wb_cpu_rdt[26] ;
 wire \u_arbiter.i_wb_cpu_rdt[27] ;
 wire \u_arbiter.i_wb_cpu_rdt[28] ;
 wire \u_arbiter.i_wb_cpu_rdt[29] ;
 wire \u_arbiter.i_wb_cpu_rdt[2] ;
 wire \u_arbiter.i_wb_cpu_rdt[30] ;
 wire \u_arbiter.i_wb_cpu_rdt[31] ;
 wire \u_arbiter.i_wb_cpu_rdt[3] ;
 wire \u_arbiter.i_wb_cpu_rdt[4] ;
 wire \u_arbiter.i_wb_cpu_rdt[5] ;
 wire \u_arbiter.i_wb_cpu_rdt[6] ;
 wire \u_arbiter.i_wb_cpu_rdt[7] ;
 wire \u_arbiter.i_wb_cpu_rdt[8] ;
 wire \u_arbiter.i_wb_cpu_rdt[9] ;
 wire \u_cpu.cpu.alu.add_cy_r ;
 wire \u_cpu.cpu.alu.cmp_r ;
 wire \u_cpu.cpu.alu.i_rs1 ;
 wire \u_cpu.cpu.bne_or_bge ;
 wire \u_cpu.cpu.branch_op ;
 wire \u_cpu.cpu.bufreg.c_r ;
 wire \u_cpu.cpu.bufreg.i_sh_signed ;
 wire \u_cpu.cpu.bufreg.lsb[0] ;
 wire \u_cpu.cpu.bufreg.lsb[1] ;
 wire \u_cpu.cpu.bufreg2.i_cnt_done ;
 wire \u_cpu.cpu.csr_d_sel ;
 wire \u_cpu.cpu.csr_imm ;
 wire \u_cpu.cpu.ctrl.i_iscomp ;
 wire \u_cpu.cpu.ctrl.i_jump ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[10] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[11] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[12] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[13] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[14] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[15] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[16] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[17] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[18] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[19] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[20] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[21] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[22] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[23] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[24] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[25] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[26] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[27] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[28] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[29] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[2] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[30] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[31] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[3] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[4] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[5] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[6] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[7] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[8] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[9] ;
 wire \u_cpu.cpu.ctrl.pc_plus_4_cy_r ;
 wire \u_cpu.cpu.ctrl.pc_plus_offset_cy_r ;
 wire \u_cpu.cpu.decode.co_ebreak ;
 wire \u_cpu.cpu.decode.co_mem_word ;
 wire \u_cpu.cpu.decode.op21 ;
 wire \u_cpu.cpu.decode.op22 ;
 wire \u_cpu.cpu.decode.op26 ;
 wire \u_cpu.cpu.decode.opcode[0] ;
 wire \u_cpu.cpu.decode.opcode[1] ;
 wire \u_cpu.cpu.decode.opcode[2] ;
 wire \u_cpu.cpu.genblk1.align.ctrl_misal ;
 wire \u_cpu.cpu.genblk1.align.ibus_rdt_concat[0] ;
 wire \u_cpu.cpu.genblk1.align.ibus_rdt_concat[10] ;
 wire \u_cpu.cpu.genblk1.align.ibus_rdt_concat[11] ;
 wire \u_cpu.cpu.genblk1.align.ibus_rdt_concat[12] ;
 wire \u_cpu.cpu.genblk1.align.ibus_rdt_concat[13] ;
 wire \u_cpu.cpu.genblk1.align.ibus_rdt_concat[14] ;
 wire \u_cpu.cpu.genblk1.align.ibus_rdt_concat[15] ;
 wire \u_cpu.cpu.genblk1.align.ibus_rdt_concat[1] ;
 wire \u_cpu.cpu.genblk1.align.ibus_rdt_concat[2] ;
 wire \u_cpu.cpu.genblk1.align.ibus_rdt_concat[3] ;
 wire \u_cpu.cpu.genblk1.align.ibus_rdt_concat[4] ;
 wire \u_cpu.cpu.genblk1.align.ibus_rdt_concat[5] ;
 wire \u_cpu.cpu.genblk1.align.ibus_rdt_concat[6] ;
 wire \u_cpu.cpu.genblk1.align.ibus_rdt_concat[7] ;
 wire \u_cpu.cpu.genblk1.align.ibus_rdt_concat[8] ;
 wire \u_cpu.cpu.genblk1.align.ibus_rdt_concat[9] ;
 wire \u_cpu.cpu.genblk3.csr.i_mtip ;
 wire \u_cpu.cpu.genblk3.csr.mcause31 ;
 wire \u_cpu.cpu.genblk3.csr.mcause3_0[0] ;
 wire \u_cpu.cpu.genblk3.csr.mcause3_0[1] ;
 wire \u_cpu.cpu.genblk3.csr.mcause3_0[2] ;
 wire \u_cpu.cpu.genblk3.csr.mcause3_0[3] ;
 wire \u_cpu.cpu.genblk3.csr.mie_mtie ;
 wire \u_cpu.cpu.genblk3.csr.mstatus_mie ;
 wire \u_cpu.cpu.genblk3.csr.mstatus_mpie ;
 wire \u_cpu.cpu.genblk3.csr.o_new_irq ;
 wire \u_cpu.cpu.genblk3.csr.timer_irq_r ;
 wire \u_cpu.cpu.immdec.imm11_7[0] ;
 wire \u_cpu.cpu.immdec.imm11_7[1] ;
 wire \u_cpu.cpu.immdec.imm11_7[2] ;
 wire \u_cpu.cpu.immdec.imm11_7[3] ;
 wire \u_cpu.cpu.immdec.imm11_7[4] ;
 wire \u_cpu.cpu.immdec.imm19_12_20[0] ;
 wire \u_cpu.cpu.immdec.imm19_12_20[1] ;
 wire \u_cpu.cpu.immdec.imm19_12_20[2] ;
 wire \u_cpu.cpu.immdec.imm19_12_20[3] ;
 wire \u_cpu.cpu.immdec.imm19_12_20[5] ;
 wire \u_cpu.cpu.immdec.imm19_12_20[6] ;
 wire \u_cpu.cpu.immdec.imm19_12_20[7] ;
 wire \u_cpu.cpu.immdec.imm19_12_20[8] ;
 wire \u_cpu.cpu.immdec.imm24_20[0] ;
 wire \u_cpu.cpu.immdec.imm24_20[1] ;
 wire \u_cpu.cpu.immdec.imm24_20[2] ;
 wire \u_cpu.cpu.immdec.imm24_20[3] ;
 wire \u_cpu.cpu.immdec.imm24_20[4] ;
 wire \u_cpu.cpu.immdec.imm30_25[0] ;
 wire \u_cpu.cpu.immdec.imm30_25[1] ;
 wire \u_cpu.cpu.immdec.imm30_25[2] ;
 wire \u_cpu.cpu.immdec.imm30_25[3] ;
 wire \u_cpu.cpu.immdec.imm30_25[4] ;
 wire \u_cpu.cpu.immdec.imm30_25[5] ;
 wire \u_cpu.cpu.immdec.imm31 ;
 wire \u_cpu.cpu.immdec.imm7 ;
 wire \u_cpu.cpu.mem_bytecnt[0] ;
 wire \u_cpu.cpu.mem_bytecnt[1] ;
 wire \u_cpu.cpu.mem_if.signbit ;
 wire \u_cpu.cpu.o_wdata0 ;
 wire \u_cpu.cpu.o_wdata1 ;
 wire \u_cpu.cpu.o_wen0 ;
 wire \u_cpu.cpu.o_wen1 ;
 wire \u_cpu.cpu.state.genblk1.misalign_trap_sync_r ;
 wire \u_cpu.cpu.state.ibus_cyc ;
 wire \u_cpu.cpu.state.init_done ;
 wire \u_cpu.cpu.state.o_cnt[2] ;
 wire \u_cpu.cpu.state.o_cnt_r[0] ;
 wire \u_cpu.cpu.state.o_cnt_r[1] ;
 wire \u_cpu.cpu.state.o_cnt_r[2] ;
 wire \u_cpu.cpu.state.o_cnt_r[3] ;
 wire \u_cpu.cpu.state.stage_two_req ;
 wire \u_cpu.raddr[0] ;
 wire \u_cpu.raddr[1] ;
 wire \u_cpu.rf_ram.memory[0][0] ;
 wire \u_cpu.rf_ram.memory[0][1] ;
 wire \u_cpu.rf_ram.memory[0][2] ;
 wire \u_cpu.rf_ram.memory[0][3] ;
 wire \u_cpu.rf_ram.memory[0][4] ;
 wire \u_cpu.rf_ram.memory[0][5] ;
 wire \u_cpu.rf_ram.memory[0][6] ;
 wire \u_cpu.rf_ram.memory[0][7] ;
 wire \u_cpu.rf_ram.memory[100][0] ;
 wire \u_cpu.rf_ram.memory[100][1] ;
 wire \u_cpu.rf_ram.memory[100][2] ;
 wire \u_cpu.rf_ram.memory[100][3] ;
 wire \u_cpu.rf_ram.memory[100][4] ;
 wire \u_cpu.rf_ram.memory[100][5] ;
 wire \u_cpu.rf_ram.memory[100][6] ;
 wire \u_cpu.rf_ram.memory[100][7] ;
 wire \u_cpu.rf_ram.memory[101][0] ;
 wire \u_cpu.rf_ram.memory[101][1] ;
 wire \u_cpu.rf_ram.memory[101][2] ;
 wire \u_cpu.rf_ram.memory[101][3] ;
 wire \u_cpu.rf_ram.memory[101][4] ;
 wire \u_cpu.rf_ram.memory[101][5] ;
 wire \u_cpu.rf_ram.memory[101][6] ;
 wire \u_cpu.rf_ram.memory[101][7] ;
 wire \u_cpu.rf_ram.memory[102][0] ;
 wire \u_cpu.rf_ram.memory[102][1] ;
 wire \u_cpu.rf_ram.memory[102][2] ;
 wire \u_cpu.rf_ram.memory[102][3] ;
 wire \u_cpu.rf_ram.memory[102][4] ;
 wire \u_cpu.rf_ram.memory[102][5] ;
 wire \u_cpu.rf_ram.memory[102][6] ;
 wire \u_cpu.rf_ram.memory[102][7] ;
 wire \u_cpu.rf_ram.memory[103][0] ;
 wire \u_cpu.rf_ram.memory[103][1] ;
 wire \u_cpu.rf_ram.memory[103][2] ;
 wire \u_cpu.rf_ram.memory[103][3] ;
 wire \u_cpu.rf_ram.memory[103][4] ;
 wire \u_cpu.rf_ram.memory[103][5] ;
 wire \u_cpu.rf_ram.memory[103][6] ;
 wire \u_cpu.rf_ram.memory[103][7] ;
 wire \u_cpu.rf_ram.memory[104][0] ;
 wire \u_cpu.rf_ram.memory[104][1] ;
 wire \u_cpu.rf_ram.memory[104][2] ;
 wire \u_cpu.rf_ram.memory[104][3] ;
 wire \u_cpu.rf_ram.memory[104][4] ;
 wire \u_cpu.rf_ram.memory[104][5] ;
 wire \u_cpu.rf_ram.memory[104][6] ;
 wire \u_cpu.rf_ram.memory[104][7] ;
 wire \u_cpu.rf_ram.memory[105][0] ;
 wire \u_cpu.rf_ram.memory[105][1] ;
 wire \u_cpu.rf_ram.memory[105][2] ;
 wire \u_cpu.rf_ram.memory[105][3] ;
 wire \u_cpu.rf_ram.memory[105][4] ;
 wire \u_cpu.rf_ram.memory[105][5] ;
 wire \u_cpu.rf_ram.memory[105][6] ;
 wire \u_cpu.rf_ram.memory[105][7] ;
 wire \u_cpu.rf_ram.memory[106][0] ;
 wire \u_cpu.rf_ram.memory[106][1] ;
 wire \u_cpu.rf_ram.memory[106][2] ;
 wire \u_cpu.rf_ram.memory[106][3] ;
 wire \u_cpu.rf_ram.memory[106][4] ;
 wire \u_cpu.rf_ram.memory[106][5] ;
 wire \u_cpu.rf_ram.memory[106][6] ;
 wire \u_cpu.rf_ram.memory[106][7] ;
 wire \u_cpu.rf_ram.memory[107][0] ;
 wire \u_cpu.rf_ram.memory[107][1] ;
 wire \u_cpu.rf_ram.memory[107][2] ;
 wire \u_cpu.rf_ram.memory[107][3] ;
 wire \u_cpu.rf_ram.memory[107][4] ;
 wire \u_cpu.rf_ram.memory[107][5] ;
 wire \u_cpu.rf_ram.memory[107][6] ;
 wire \u_cpu.rf_ram.memory[107][7] ;
 wire \u_cpu.rf_ram.memory[108][0] ;
 wire \u_cpu.rf_ram.memory[108][1] ;
 wire \u_cpu.rf_ram.memory[108][2] ;
 wire \u_cpu.rf_ram.memory[108][3] ;
 wire \u_cpu.rf_ram.memory[108][4] ;
 wire \u_cpu.rf_ram.memory[108][5] ;
 wire \u_cpu.rf_ram.memory[108][6] ;
 wire \u_cpu.rf_ram.memory[108][7] ;
 wire \u_cpu.rf_ram.memory[109][0] ;
 wire \u_cpu.rf_ram.memory[109][1] ;
 wire \u_cpu.rf_ram.memory[109][2] ;
 wire \u_cpu.rf_ram.memory[109][3] ;
 wire \u_cpu.rf_ram.memory[109][4] ;
 wire \u_cpu.rf_ram.memory[109][5] ;
 wire \u_cpu.rf_ram.memory[109][6] ;
 wire \u_cpu.rf_ram.memory[109][7] ;
 wire \u_cpu.rf_ram.memory[10][0] ;
 wire \u_cpu.rf_ram.memory[10][1] ;
 wire \u_cpu.rf_ram.memory[10][2] ;
 wire \u_cpu.rf_ram.memory[10][3] ;
 wire \u_cpu.rf_ram.memory[10][4] ;
 wire \u_cpu.rf_ram.memory[10][5] ;
 wire \u_cpu.rf_ram.memory[10][6] ;
 wire \u_cpu.rf_ram.memory[10][7] ;
 wire \u_cpu.rf_ram.memory[110][0] ;
 wire \u_cpu.rf_ram.memory[110][1] ;
 wire \u_cpu.rf_ram.memory[110][2] ;
 wire \u_cpu.rf_ram.memory[110][3] ;
 wire \u_cpu.rf_ram.memory[110][4] ;
 wire \u_cpu.rf_ram.memory[110][5] ;
 wire \u_cpu.rf_ram.memory[110][6] ;
 wire \u_cpu.rf_ram.memory[110][7] ;
 wire \u_cpu.rf_ram.memory[111][0] ;
 wire \u_cpu.rf_ram.memory[111][1] ;
 wire \u_cpu.rf_ram.memory[111][2] ;
 wire \u_cpu.rf_ram.memory[111][3] ;
 wire \u_cpu.rf_ram.memory[111][4] ;
 wire \u_cpu.rf_ram.memory[111][5] ;
 wire \u_cpu.rf_ram.memory[111][6] ;
 wire \u_cpu.rf_ram.memory[111][7] ;
 wire \u_cpu.rf_ram.memory[112][0] ;
 wire \u_cpu.rf_ram.memory[112][1] ;
 wire \u_cpu.rf_ram.memory[112][2] ;
 wire \u_cpu.rf_ram.memory[112][3] ;
 wire \u_cpu.rf_ram.memory[112][4] ;
 wire \u_cpu.rf_ram.memory[112][5] ;
 wire \u_cpu.rf_ram.memory[112][6] ;
 wire \u_cpu.rf_ram.memory[112][7] ;
 wire \u_cpu.rf_ram.memory[113][0] ;
 wire \u_cpu.rf_ram.memory[113][1] ;
 wire \u_cpu.rf_ram.memory[113][2] ;
 wire \u_cpu.rf_ram.memory[113][3] ;
 wire \u_cpu.rf_ram.memory[113][4] ;
 wire \u_cpu.rf_ram.memory[113][5] ;
 wire \u_cpu.rf_ram.memory[113][6] ;
 wire \u_cpu.rf_ram.memory[113][7] ;
 wire \u_cpu.rf_ram.memory[114][0] ;
 wire \u_cpu.rf_ram.memory[114][1] ;
 wire \u_cpu.rf_ram.memory[114][2] ;
 wire \u_cpu.rf_ram.memory[114][3] ;
 wire \u_cpu.rf_ram.memory[114][4] ;
 wire \u_cpu.rf_ram.memory[114][5] ;
 wire \u_cpu.rf_ram.memory[114][6] ;
 wire \u_cpu.rf_ram.memory[114][7] ;
 wire \u_cpu.rf_ram.memory[115][0] ;
 wire \u_cpu.rf_ram.memory[115][1] ;
 wire \u_cpu.rf_ram.memory[115][2] ;
 wire \u_cpu.rf_ram.memory[115][3] ;
 wire \u_cpu.rf_ram.memory[115][4] ;
 wire \u_cpu.rf_ram.memory[115][5] ;
 wire \u_cpu.rf_ram.memory[115][6] ;
 wire \u_cpu.rf_ram.memory[115][7] ;
 wire \u_cpu.rf_ram.memory[116][0] ;
 wire \u_cpu.rf_ram.memory[116][1] ;
 wire \u_cpu.rf_ram.memory[116][2] ;
 wire \u_cpu.rf_ram.memory[116][3] ;
 wire \u_cpu.rf_ram.memory[116][4] ;
 wire \u_cpu.rf_ram.memory[116][5] ;
 wire \u_cpu.rf_ram.memory[116][6] ;
 wire \u_cpu.rf_ram.memory[116][7] ;
 wire \u_cpu.rf_ram.memory[117][0] ;
 wire \u_cpu.rf_ram.memory[117][1] ;
 wire \u_cpu.rf_ram.memory[117][2] ;
 wire \u_cpu.rf_ram.memory[117][3] ;
 wire \u_cpu.rf_ram.memory[117][4] ;
 wire \u_cpu.rf_ram.memory[117][5] ;
 wire \u_cpu.rf_ram.memory[117][6] ;
 wire \u_cpu.rf_ram.memory[117][7] ;
 wire \u_cpu.rf_ram.memory[118][0] ;
 wire \u_cpu.rf_ram.memory[118][1] ;
 wire \u_cpu.rf_ram.memory[118][2] ;
 wire \u_cpu.rf_ram.memory[118][3] ;
 wire \u_cpu.rf_ram.memory[118][4] ;
 wire \u_cpu.rf_ram.memory[118][5] ;
 wire \u_cpu.rf_ram.memory[118][6] ;
 wire \u_cpu.rf_ram.memory[118][7] ;
 wire \u_cpu.rf_ram.memory[119][0] ;
 wire \u_cpu.rf_ram.memory[119][1] ;
 wire \u_cpu.rf_ram.memory[119][2] ;
 wire \u_cpu.rf_ram.memory[119][3] ;
 wire \u_cpu.rf_ram.memory[119][4] ;
 wire \u_cpu.rf_ram.memory[119][5] ;
 wire \u_cpu.rf_ram.memory[119][6] ;
 wire \u_cpu.rf_ram.memory[119][7] ;
 wire \u_cpu.rf_ram.memory[11][0] ;
 wire \u_cpu.rf_ram.memory[11][1] ;
 wire \u_cpu.rf_ram.memory[11][2] ;
 wire \u_cpu.rf_ram.memory[11][3] ;
 wire \u_cpu.rf_ram.memory[11][4] ;
 wire \u_cpu.rf_ram.memory[11][5] ;
 wire \u_cpu.rf_ram.memory[11][6] ;
 wire \u_cpu.rf_ram.memory[11][7] ;
 wire \u_cpu.rf_ram.memory[120][0] ;
 wire \u_cpu.rf_ram.memory[120][1] ;
 wire \u_cpu.rf_ram.memory[120][2] ;
 wire \u_cpu.rf_ram.memory[120][3] ;
 wire \u_cpu.rf_ram.memory[120][4] ;
 wire \u_cpu.rf_ram.memory[120][5] ;
 wire \u_cpu.rf_ram.memory[120][6] ;
 wire \u_cpu.rf_ram.memory[120][7] ;
 wire \u_cpu.rf_ram.memory[121][0] ;
 wire \u_cpu.rf_ram.memory[121][1] ;
 wire \u_cpu.rf_ram.memory[121][2] ;
 wire \u_cpu.rf_ram.memory[121][3] ;
 wire \u_cpu.rf_ram.memory[121][4] ;
 wire \u_cpu.rf_ram.memory[121][5] ;
 wire \u_cpu.rf_ram.memory[121][6] ;
 wire \u_cpu.rf_ram.memory[121][7] ;
 wire \u_cpu.rf_ram.memory[122][0] ;
 wire \u_cpu.rf_ram.memory[122][1] ;
 wire \u_cpu.rf_ram.memory[122][2] ;
 wire \u_cpu.rf_ram.memory[122][3] ;
 wire \u_cpu.rf_ram.memory[122][4] ;
 wire \u_cpu.rf_ram.memory[122][5] ;
 wire \u_cpu.rf_ram.memory[122][6] ;
 wire \u_cpu.rf_ram.memory[122][7] ;
 wire \u_cpu.rf_ram.memory[123][0] ;
 wire \u_cpu.rf_ram.memory[123][1] ;
 wire \u_cpu.rf_ram.memory[123][2] ;
 wire \u_cpu.rf_ram.memory[123][3] ;
 wire \u_cpu.rf_ram.memory[123][4] ;
 wire \u_cpu.rf_ram.memory[123][5] ;
 wire \u_cpu.rf_ram.memory[123][6] ;
 wire \u_cpu.rf_ram.memory[123][7] ;
 wire \u_cpu.rf_ram.memory[124][0] ;
 wire \u_cpu.rf_ram.memory[124][1] ;
 wire \u_cpu.rf_ram.memory[124][2] ;
 wire \u_cpu.rf_ram.memory[124][3] ;
 wire \u_cpu.rf_ram.memory[124][4] ;
 wire \u_cpu.rf_ram.memory[124][5] ;
 wire \u_cpu.rf_ram.memory[124][6] ;
 wire \u_cpu.rf_ram.memory[124][7] ;
 wire \u_cpu.rf_ram.memory[125][0] ;
 wire \u_cpu.rf_ram.memory[125][1] ;
 wire \u_cpu.rf_ram.memory[125][2] ;
 wire \u_cpu.rf_ram.memory[125][3] ;
 wire \u_cpu.rf_ram.memory[125][4] ;
 wire \u_cpu.rf_ram.memory[125][5] ;
 wire \u_cpu.rf_ram.memory[125][6] ;
 wire \u_cpu.rf_ram.memory[125][7] ;
 wire \u_cpu.rf_ram.memory[126][0] ;
 wire \u_cpu.rf_ram.memory[126][1] ;
 wire \u_cpu.rf_ram.memory[126][2] ;
 wire \u_cpu.rf_ram.memory[126][3] ;
 wire \u_cpu.rf_ram.memory[126][4] ;
 wire \u_cpu.rf_ram.memory[126][5] ;
 wire \u_cpu.rf_ram.memory[126][6] ;
 wire \u_cpu.rf_ram.memory[126][7] ;
 wire \u_cpu.rf_ram.memory[127][0] ;
 wire \u_cpu.rf_ram.memory[127][1] ;
 wire \u_cpu.rf_ram.memory[127][2] ;
 wire \u_cpu.rf_ram.memory[127][3] ;
 wire \u_cpu.rf_ram.memory[127][4] ;
 wire \u_cpu.rf_ram.memory[127][5] ;
 wire \u_cpu.rf_ram.memory[127][6] ;
 wire \u_cpu.rf_ram.memory[127][7] ;
 wire \u_cpu.rf_ram.memory[128][0] ;
 wire \u_cpu.rf_ram.memory[128][1] ;
 wire \u_cpu.rf_ram.memory[128][2] ;
 wire \u_cpu.rf_ram.memory[128][3] ;
 wire \u_cpu.rf_ram.memory[128][4] ;
 wire \u_cpu.rf_ram.memory[128][5] ;
 wire \u_cpu.rf_ram.memory[128][6] ;
 wire \u_cpu.rf_ram.memory[128][7] ;
 wire \u_cpu.rf_ram.memory[129][0] ;
 wire \u_cpu.rf_ram.memory[129][1] ;
 wire \u_cpu.rf_ram.memory[129][2] ;
 wire \u_cpu.rf_ram.memory[129][3] ;
 wire \u_cpu.rf_ram.memory[129][4] ;
 wire \u_cpu.rf_ram.memory[129][5] ;
 wire \u_cpu.rf_ram.memory[129][6] ;
 wire \u_cpu.rf_ram.memory[129][7] ;
 wire \u_cpu.rf_ram.memory[12][0] ;
 wire \u_cpu.rf_ram.memory[12][1] ;
 wire \u_cpu.rf_ram.memory[12][2] ;
 wire \u_cpu.rf_ram.memory[12][3] ;
 wire \u_cpu.rf_ram.memory[12][4] ;
 wire \u_cpu.rf_ram.memory[12][5] ;
 wire \u_cpu.rf_ram.memory[12][6] ;
 wire \u_cpu.rf_ram.memory[12][7] ;
 wire \u_cpu.rf_ram.memory[130][0] ;
 wire \u_cpu.rf_ram.memory[130][1] ;
 wire \u_cpu.rf_ram.memory[130][2] ;
 wire \u_cpu.rf_ram.memory[130][3] ;
 wire \u_cpu.rf_ram.memory[130][4] ;
 wire \u_cpu.rf_ram.memory[130][5] ;
 wire \u_cpu.rf_ram.memory[130][6] ;
 wire \u_cpu.rf_ram.memory[130][7] ;
 wire \u_cpu.rf_ram.memory[131][0] ;
 wire \u_cpu.rf_ram.memory[131][1] ;
 wire \u_cpu.rf_ram.memory[131][2] ;
 wire \u_cpu.rf_ram.memory[131][3] ;
 wire \u_cpu.rf_ram.memory[131][4] ;
 wire \u_cpu.rf_ram.memory[131][5] ;
 wire \u_cpu.rf_ram.memory[131][6] ;
 wire \u_cpu.rf_ram.memory[131][7] ;
 wire \u_cpu.rf_ram.memory[132][0] ;
 wire \u_cpu.rf_ram.memory[132][1] ;
 wire \u_cpu.rf_ram.memory[132][2] ;
 wire \u_cpu.rf_ram.memory[132][3] ;
 wire \u_cpu.rf_ram.memory[132][4] ;
 wire \u_cpu.rf_ram.memory[132][5] ;
 wire \u_cpu.rf_ram.memory[132][6] ;
 wire \u_cpu.rf_ram.memory[132][7] ;
 wire \u_cpu.rf_ram.memory[133][0] ;
 wire \u_cpu.rf_ram.memory[133][1] ;
 wire \u_cpu.rf_ram.memory[133][2] ;
 wire \u_cpu.rf_ram.memory[133][3] ;
 wire \u_cpu.rf_ram.memory[133][4] ;
 wire \u_cpu.rf_ram.memory[133][5] ;
 wire \u_cpu.rf_ram.memory[133][6] ;
 wire \u_cpu.rf_ram.memory[133][7] ;
 wire \u_cpu.rf_ram.memory[134][0] ;
 wire \u_cpu.rf_ram.memory[134][1] ;
 wire \u_cpu.rf_ram.memory[134][2] ;
 wire \u_cpu.rf_ram.memory[134][3] ;
 wire \u_cpu.rf_ram.memory[134][4] ;
 wire \u_cpu.rf_ram.memory[134][5] ;
 wire \u_cpu.rf_ram.memory[134][6] ;
 wire \u_cpu.rf_ram.memory[134][7] ;
 wire \u_cpu.rf_ram.memory[135][0] ;
 wire \u_cpu.rf_ram.memory[135][1] ;
 wire \u_cpu.rf_ram.memory[135][2] ;
 wire \u_cpu.rf_ram.memory[135][3] ;
 wire \u_cpu.rf_ram.memory[135][4] ;
 wire \u_cpu.rf_ram.memory[135][5] ;
 wire \u_cpu.rf_ram.memory[135][6] ;
 wire \u_cpu.rf_ram.memory[135][7] ;
 wire \u_cpu.rf_ram.memory[136][0] ;
 wire \u_cpu.rf_ram.memory[136][1] ;
 wire \u_cpu.rf_ram.memory[136][2] ;
 wire \u_cpu.rf_ram.memory[136][3] ;
 wire \u_cpu.rf_ram.memory[136][4] ;
 wire \u_cpu.rf_ram.memory[136][5] ;
 wire \u_cpu.rf_ram.memory[136][6] ;
 wire \u_cpu.rf_ram.memory[136][7] ;
 wire \u_cpu.rf_ram.memory[137][0] ;
 wire \u_cpu.rf_ram.memory[137][1] ;
 wire \u_cpu.rf_ram.memory[137][2] ;
 wire \u_cpu.rf_ram.memory[137][3] ;
 wire \u_cpu.rf_ram.memory[137][4] ;
 wire \u_cpu.rf_ram.memory[137][5] ;
 wire \u_cpu.rf_ram.memory[137][6] ;
 wire \u_cpu.rf_ram.memory[137][7] ;
 wire \u_cpu.rf_ram.memory[138][0] ;
 wire \u_cpu.rf_ram.memory[138][1] ;
 wire \u_cpu.rf_ram.memory[138][2] ;
 wire \u_cpu.rf_ram.memory[138][3] ;
 wire \u_cpu.rf_ram.memory[138][4] ;
 wire \u_cpu.rf_ram.memory[138][5] ;
 wire \u_cpu.rf_ram.memory[138][6] ;
 wire \u_cpu.rf_ram.memory[138][7] ;
 wire \u_cpu.rf_ram.memory[139][0] ;
 wire \u_cpu.rf_ram.memory[139][1] ;
 wire \u_cpu.rf_ram.memory[139][2] ;
 wire \u_cpu.rf_ram.memory[139][3] ;
 wire \u_cpu.rf_ram.memory[139][4] ;
 wire \u_cpu.rf_ram.memory[139][5] ;
 wire \u_cpu.rf_ram.memory[139][6] ;
 wire \u_cpu.rf_ram.memory[139][7] ;
 wire \u_cpu.rf_ram.memory[13][0] ;
 wire \u_cpu.rf_ram.memory[13][1] ;
 wire \u_cpu.rf_ram.memory[13][2] ;
 wire \u_cpu.rf_ram.memory[13][3] ;
 wire \u_cpu.rf_ram.memory[13][4] ;
 wire \u_cpu.rf_ram.memory[13][5] ;
 wire \u_cpu.rf_ram.memory[13][6] ;
 wire \u_cpu.rf_ram.memory[13][7] ;
 wire \u_cpu.rf_ram.memory[140][0] ;
 wire \u_cpu.rf_ram.memory[140][1] ;
 wire \u_cpu.rf_ram.memory[140][2] ;
 wire \u_cpu.rf_ram.memory[140][3] ;
 wire \u_cpu.rf_ram.memory[140][4] ;
 wire \u_cpu.rf_ram.memory[140][5] ;
 wire \u_cpu.rf_ram.memory[140][6] ;
 wire \u_cpu.rf_ram.memory[140][7] ;
 wire \u_cpu.rf_ram.memory[141][0] ;
 wire \u_cpu.rf_ram.memory[141][1] ;
 wire \u_cpu.rf_ram.memory[141][2] ;
 wire \u_cpu.rf_ram.memory[141][3] ;
 wire \u_cpu.rf_ram.memory[141][4] ;
 wire \u_cpu.rf_ram.memory[141][5] ;
 wire \u_cpu.rf_ram.memory[141][6] ;
 wire \u_cpu.rf_ram.memory[141][7] ;
 wire \u_cpu.rf_ram.memory[142][0] ;
 wire \u_cpu.rf_ram.memory[142][1] ;
 wire \u_cpu.rf_ram.memory[142][2] ;
 wire \u_cpu.rf_ram.memory[142][3] ;
 wire \u_cpu.rf_ram.memory[142][4] ;
 wire \u_cpu.rf_ram.memory[142][5] ;
 wire \u_cpu.rf_ram.memory[142][6] ;
 wire \u_cpu.rf_ram.memory[142][7] ;
 wire \u_cpu.rf_ram.memory[143][0] ;
 wire \u_cpu.rf_ram.memory[143][1] ;
 wire \u_cpu.rf_ram.memory[143][2] ;
 wire \u_cpu.rf_ram.memory[143][3] ;
 wire \u_cpu.rf_ram.memory[143][4] ;
 wire \u_cpu.rf_ram.memory[143][5] ;
 wire \u_cpu.rf_ram.memory[143][6] ;
 wire \u_cpu.rf_ram.memory[143][7] ;
 wire \u_cpu.rf_ram.memory[14][0] ;
 wire \u_cpu.rf_ram.memory[14][1] ;
 wire \u_cpu.rf_ram.memory[14][2] ;
 wire \u_cpu.rf_ram.memory[14][3] ;
 wire \u_cpu.rf_ram.memory[14][4] ;
 wire \u_cpu.rf_ram.memory[14][5] ;
 wire \u_cpu.rf_ram.memory[14][6] ;
 wire \u_cpu.rf_ram.memory[14][7] ;
 wire \u_cpu.rf_ram.memory[15][0] ;
 wire \u_cpu.rf_ram.memory[15][1] ;
 wire \u_cpu.rf_ram.memory[15][2] ;
 wire \u_cpu.rf_ram.memory[15][3] ;
 wire \u_cpu.rf_ram.memory[15][4] ;
 wire \u_cpu.rf_ram.memory[15][5] ;
 wire \u_cpu.rf_ram.memory[15][6] ;
 wire \u_cpu.rf_ram.memory[15][7] ;
 wire \u_cpu.rf_ram.memory[16][0] ;
 wire \u_cpu.rf_ram.memory[16][1] ;
 wire \u_cpu.rf_ram.memory[16][2] ;
 wire \u_cpu.rf_ram.memory[16][3] ;
 wire \u_cpu.rf_ram.memory[16][4] ;
 wire \u_cpu.rf_ram.memory[16][5] ;
 wire \u_cpu.rf_ram.memory[16][6] ;
 wire \u_cpu.rf_ram.memory[16][7] ;
 wire \u_cpu.rf_ram.memory[17][0] ;
 wire \u_cpu.rf_ram.memory[17][1] ;
 wire \u_cpu.rf_ram.memory[17][2] ;
 wire \u_cpu.rf_ram.memory[17][3] ;
 wire \u_cpu.rf_ram.memory[17][4] ;
 wire \u_cpu.rf_ram.memory[17][5] ;
 wire \u_cpu.rf_ram.memory[17][6] ;
 wire \u_cpu.rf_ram.memory[17][7] ;
 wire \u_cpu.rf_ram.memory[18][0] ;
 wire \u_cpu.rf_ram.memory[18][1] ;
 wire \u_cpu.rf_ram.memory[18][2] ;
 wire \u_cpu.rf_ram.memory[18][3] ;
 wire \u_cpu.rf_ram.memory[18][4] ;
 wire \u_cpu.rf_ram.memory[18][5] ;
 wire \u_cpu.rf_ram.memory[18][6] ;
 wire \u_cpu.rf_ram.memory[18][7] ;
 wire \u_cpu.rf_ram.memory[19][0] ;
 wire \u_cpu.rf_ram.memory[19][1] ;
 wire \u_cpu.rf_ram.memory[19][2] ;
 wire \u_cpu.rf_ram.memory[19][3] ;
 wire \u_cpu.rf_ram.memory[19][4] ;
 wire \u_cpu.rf_ram.memory[19][5] ;
 wire \u_cpu.rf_ram.memory[19][6] ;
 wire \u_cpu.rf_ram.memory[19][7] ;
 wire \u_cpu.rf_ram.memory[1][0] ;
 wire \u_cpu.rf_ram.memory[1][1] ;
 wire \u_cpu.rf_ram.memory[1][2] ;
 wire \u_cpu.rf_ram.memory[1][3] ;
 wire \u_cpu.rf_ram.memory[1][4] ;
 wire \u_cpu.rf_ram.memory[1][5] ;
 wire \u_cpu.rf_ram.memory[1][6] ;
 wire \u_cpu.rf_ram.memory[1][7] ;
 wire \u_cpu.rf_ram.memory[20][0] ;
 wire \u_cpu.rf_ram.memory[20][1] ;
 wire \u_cpu.rf_ram.memory[20][2] ;
 wire \u_cpu.rf_ram.memory[20][3] ;
 wire \u_cpu.rf_ram.memory[20][4] ;
 wire \u_cpu.rf_ram.memory[20][5] ;
 wire \u_cpu.rf_ram.memory[20][6] ;
 wire \u_cpu.rf_ram.memory[20][7] ;
 wire \u_cpu.rf_ram.memory[21][0] ;
 wire \u_cpu.rf_ram.memory[21][1] ;
 wire \u_cpu.rf_ram.memory[21][2] ;
 wire \u_cpu.rf_ram.memory[21][3] ;
 wire \u_cpu.rf_ram.memory[21][4] ;
 wire \u_cpu.rf_ram.memory[21][5] ;
 wire \u_cpu.rf_ram.memory[21][6] ;
 wire \u_cpu.rf_ram.memory[21][7] ;
 wire \u_cpu.rf_ram.memory[22][0] ;
 wire \u_cpu.rf_ram.memory[22][1] ;
 wire \u_cpu.rf_ram.memory[22][2] ;
 wire \u_cpu.rf_ram.memory[22][3] ;
 wire \u_cpu.rf_ram.memory[22][4] ;
 wire \u_cpu.rf_ram.memory[22][5] ;
 wire \u_cpu.rf_ram.memory[22][6] ;
 wire \u_cpu.rf_ram.memory[22][7] ;
 wire \u_cpu.rf_ram.memory[23][0] ;
 wire \u_cpu.rf_ram.memory[23][1] ;
 wire \u_cpu.rf_ram.memory[23][2] ;
 wire \u_cpu.rf_ram.memory[23][3] ;
 wire \u_cpu.rf_ram.memory[23][4] ;
 wire \u_cpu.rf_ram.memory[23][5] ;
 wire \u_cpu.rf_ram.memory[23][6] ;
 wire \u_cpu.rf_ram.memory[23][7] ;
 wire \u_cpu.rf_ram.memory[24][0] ;
 wire \u_cpu.rf_ram.memory[24][1] ;
 wire \u_cpu.rf_ram.memory[24][2] ;
 wire \u_cpu.rf_ram.memory[24][3] ;
 wire \u_cpu.rf_ram.memory[24][4] ;
 wire \u_cpu.rf_ram.memory[24][5] ;
 wire \u_cpu.rf_ram.memory[24][6] ;
 wire \u_cpu.rf_ram.memory[24][7] ;
 wire \u_cpu.rf_ram.memory[25][0] ;
 wire \u_cpu.rf_ram.memory[25][1] ;
 wire \u_cpu.rf_ram.memory[25][2] ;
 wire \u_cpu.rf_ram.memory[25][3] ;
 wire \u_cpu.rf_ram.memory[25][4] ;
 wire \u_cpu.rf_ram.memory[25][5] ;
 wire \u_cpu.rf_ram.memory[25][6] ;
 wire \u_cpu.rf_ram.memory[25][7] ;
 wire \u_cpu.rf_ram.memory[26][0] ;
 wire \u_cpu.rf_ram.memory[26][1] ;
 wire \u_cpu.rf_ram.memory[26][2] ;
 wire \u_cpu.rf_ram.memory[26][3] ;
 wire \u_cpu.rf_ram.memory[26][4] ;
 wire \u_cpu.rf_ram.memory[26][5] ;
 wire \u_cpu.rf_ram.memory[26][6] ;
 wire \u_cpu.rf_ram.memory[26][7] ;
 wire \u_cpu.rf_ram.memory[27][0] ;
 wire \u_cpu.rf_ram.memory[27][1] ;
 wire \u_cpu.rf_ram.memory[27][2] ;
 wire \u_cpu.rf_ram.memory[27][3] ;
 wire \u_cpu.rf_ram.memory[27][4] ;
 wire \u_cpu.rf_ram.memory[27][5] ;
 wire \u_cpu.rf_ram.memory[27][6] ;
 wire \u_cpu.rf_ram.memory[27][7] ;
 wire \u_cpu.rf_ram.memory[28][0] ;
 wire \u_cpu.rf_ram.memory[28][1] ;
 wire \u_cpu.rf_ram.memory[28][2] ;
 wire \u_cpu.rf_ram.memory[28][3] ;
 wire \u_cpu.rf_ram.memory[28][4] ;
 wire \u_cpu.rf_ram.memory[28][5] ;
 wire \u_cpu.rf_ram.memory[28][6] ;
 wire \u_cpu.rf_ram.memory[28][7] ;
 wire \u_cpu.rf_ram.memory[29][0] ;
 wire \u_cpu.rf_ram.memory[29][1] ;
 wire \u_cpu.rf_ram.memory[29][2] ;
 wire \u_cpu.rf_ram.memory[29][3] ;
 wire \u_cpu.rf_ram.memory[29][4] ;
 wire \u_cpu.rf_ram.memory[29][5] ;
 wire \u_cpu.rf_ram.memory[29][6] ;
 wire \u_cpu.rf_ram.memory[29][7] ;
 wire \u_cpu.rf_ram.memory[2][0] ;
 wire \u_cpu.rf_ram.memory[2][1] ;
 wire \u_cpu.rf_ram.memory[2][2] ;
 wire \u_cpu.rf_ram.memory[2][3] ;
 wire \u_cpu.rf_ram.memory[2][4] ;
 wire \u_cpu.rf_ram.memory[2][5] ;
 wire \u_cpu.rf_ram.memory[2][6] ;
 wire \u_cpu.rf_ram.memory[2][7] ;
 wire \u_cpu.rf_ram.memory[30][0] ;
 wire \u_cpu.rf_ram.memory[30][1] ;
 wire \u_cpu.rf_ram.memory[30][2] ;
 wire \u_cpu.rf_ram.memory[30][3] ;
 wire \u_cpu.rf_ram.memory[30][4] ;
 wire \u_cpu.rf_ram.memory[30][5] ;
 wire \u_cpu.rf_ram.memory[30][6] ;
 wire \u_cpu.rf_ram.memory[30][7] ;
 wire \u_cpu.rf_ram.memory[31][0] ;
 wire \u_cpu.rf_ram.memory[31][1] ;
 wire \u_cpu.rf_ram.memory[31][2] ;
 wire \u_cpu.rf_ram.memory[31][3] ;
 wire \u_cpu.rf_ram.memory[31][4] ;
 wire \u_cpu.rf_ram.memory[31][5] ;
 wire \u_cpu.rf_ram.memory[31][6] ;
 wire \u_cpu.rf_ram.memory[31][7] ;
 wire \u_cpu.rf_ram.memory[32][0] ;
 wire \u_cpu.rf_ram.memory[32][1] ;
 wire \u_cpu.rf_ram.memory[32][2] ;
 wire \u_cpu.rf_ram.memory[32][3] ;
 wire \u_cpu.rf_ram.memory[32][4] ;
 wire \u_cpu.rf_ram.memory[32][5] ;
 wire \u_cpu.rf_ram.memory[32][6] ;
 wire \u_cpu.rf_ram.memory[32][7] ;
 wire \u_cpu.rf_ram.memory[33][0] ;
 wire \u_cpu.rf_ram.memory[33][1] ;
 wire \u_cpu.rf_ram.memory[33][2] ;
 wire \u_cpu.rf_ram.memory[33][3] ;
 wire \u_cpu.rf_ram.memory[33][4] ;
 wire \u_cpu.rf_ram.memory[33][5] ;
 wire \u_cpu.rf_ram.memory[33][6] ;
 wire \u_cpu.rf_ram.memory[33][7] ;
 wire \u_cpu.rf_ram.memory[34][0] ;
 wire \u_cpu.rf_ram.memory[34][1] ;
 wire \u_cpu.rf_ram.memory[34][2] ;
 wire \u_cpu.rf_ram.memory[34][3] ;
 wire \u_cpu.rf_ram.memory[34][4] ;
 wire \u_cpu.rf_ram.memory[34][5] ;
 wire \u_cpu.rf_ram.memory[34][6] ;
 wire \u_cpu.rf_ram.memory[34][7] ;
 wire \u_cpu.rf_ram.memory[35][0] ;
 wire \u_cpu.rf_ram.memory[35][1] ;
 wire \u_cpu.rf_ram.memory[35][2] ;
 wire \u_cpu.rf_ram.memory[35][3] ;
 wire \u_cpu.rf_ram.memory[35][4] ;
 wire \u_cpu.rf_ram.memory[35][5] ;
 wire \u_cpu.rf_ram.memory[35][6] ;
 wire \u_cpu.rf_ram.memory[35][7] ;
 wire \u_cpu.rf_ram.memory[36][0] ;
 wire \u_cpu.rf_ram.memory[36][1] ;
 wire \u_cpu.rf_ram.memory[36][2] ;
 wire \u_cpu.rf_ram.memory[36][3] ;
 wire \u_cpu.rf_ram.memory[36][4] ;
 wire \u_cpu.rf_ram.memory[36][5] ;
 wire \u_cpu.rf_ram.memory[36][6] ;
 wire \u_cpu.rf_ram.memory[36][7] ;
 wire \u_cpu.rf_ram.memory[37][0] ;
 wire \u_cpu.rf_ram.memory[37][1] ;
 wire \u_cpu.rf_ram.memory[37][2] ;
 wire \u_cpu.rf_ram.memory[37][3] ;
 wire \u_cpu.rf_ram.memory[37][4] ;
 wire \u_cpu.rf_ram.memory[37][5] ;
 wire \u_cpu.rf_ram.memory[37][6] ;
 wire \u_cpu.rf_ram.memory[37][7] ;
 wire \u_cpu.rf_ram.memory[38][0] ;
 wire \u_cpu.rf_ram.memory[38][1] ;
 wire \u_cpu.rf_ram.memory[38][2] ;
 wire \u_cpu.rf_ram.memory[38][3] ;
 wire \u_cpu.rf_ram.memory[38][4] ;
 wire \u_cpu.rf_ram.memory[38][5] ;
 wire \u_cpu.rf_ram.memory[38][6] ;
 wire \u_cpu.rf_ram.memory[38][7] ;
 wire \u_cpu.rf_ram.memory[39][0] ;
 wire \u_cpu.rf_ram.memory[39][1] ;
 wire \u_cpu.rf_ram.memory[39][2] ;
 wire \u_cpu.rf_ram.memory[39][3] ;
 wire \u_cpu.rf_ram.memory[39][4] ;
 wire \u_cpu.rf_ram.memory[39][5] ;
 wire \u_cpu.rf_ram.memory[39][6] ;
 wire \u_cpu.rf_ram.memory[39][7] ;
 wire \u_cpu.rf_ram.memory[3][0] ;
 wire \u_cpu.rf_ram.memory[3][1] ;
 wire \u_cpu.rf_ram.memory[3][2] ;
 wire \u_cpu.rf_ram.memory[3][3] ;
 wire \u_cpu.rf_ram.memory[3][4] ;
 wire \u_cpu.rf_ram.memory[3][5] ;
 wire \u_cpu.rf_ram.memory[3][6] ;
 wire \u_cpu.rf_ram.memory[3][7] ;
 wire \u_cpu.rf_ram.memory[40][0] ;
 wire \u_cpu.rf_ram.memory[40][1] ;
 wire \u_cpu.rf_ram.memory[40][2] ;
 wire \u_cpu.rf_ram.memory[40][3] ;
 wire \u_cpu.rf_ram.memory[40][4] ;
 wire \u_cpu.rf_ram.memory[40][5] ;
 wire \u_cpu.rf_ram.memory[40][6] ;
 wire \u_cpu.rf_ram.memory[40][7] ;
 wire \u_cpu.rf_ram.memory[41][0] ;
 wire \u_cpu.rf_ram.memory[41][1] ;
 wire \u_cpu.rf_ram.memory[41][2] ;
 wire \u_cpu.rf_ram.memory[41][3] ;
 wire \u_cpu.rf_ram.memory[41][4] ;
 wire \u_cpu.rf_ram.memory[41][5] ;
 wire \u_cpu.rf_ram.memory[41][6] ;
 wire \u_cpu.rf_ram.memory[41][7] ;
 wire \u_cpu.rf_ram.memory[42][0] ;
 wire \u_cpu.rf_ram.memory[42][1] ;
 wire \u_cpu.rf_ram.memory[42][2] ;
 wire \u_cpu.rf_ram.memory[42][3] ;
 wire \u_cpu.rf_ram.memory[42][4] ;
 wire \u_cpu.rf_ram.memory[42][5] ;
 wire \u_cpu.rf_ram.memory[42][6] ;
 wire \u_cpu.rf_ram.memory[42][7] ;
 wire \u_cpu.rf_ram.memory[43][0] ;
 wire \u_cpu.rf_ram.memory[43][1] ;
 wire \u_cpu.rf_ram.memory[43][2] ;
 wire \u_cpu.rf_ram.memory[43][3] ;
 wire \u_cpu.rf_ram.memory[43][4] ;
 wire \u_cpu.rf_ram.memory[43][5] ;
 wire \u_cpu.rf_ram.memory[43][6] ;
 wire \u_cpu.rf_ram.memory[43][7] ;
 wire \u_cpu.rf_ram.memory[44][0] ;
 wire \u_cpu.rf_ram.memory[44][1] ;
 wire \u_cpu.rf_ram.memory[44][2] ;
 wire \u_cpu.rf_ram.memory[44][3] ;
 wire \u_cpu.rf_ram.memory[44][4] ;
 wire \u_cpu.rf_ram.memory[44][5] ;
 wire \u_cpu.rf_ram.memory[44][6] ;
 wire \u_cpu.rf_ram.memory[44][7] ;
 wire \u_cpu.rf_ram.memory[45][0] ;
 wire \u_cpu.rf_ram.memory[45][1] ;
 wire \u_cpu.rf_ram.memory[45][2] ;
 wire \u_cpu.rf_ram.memory[45][3] ;
 wire \u_cpu.rf_ram.memory[45][4] ;
 wire \u_cpu.rf_ram.memory[45][5] ;
 wire \u_cpu.rf_ram.memory[45][6] ;
 wire \u_cpu.rf_ram.memory[45][7] ;
 wire \u_cpu.rf_ram.memory[46][0] ;
 wire \u_cpu.rf_ram.memory[46][1] ;
 wire \u_cpu.rf_ram.memory[46][2] ;
 wire \u_cpu.rf_ram.memory[46][3] ;
 wire \u_cpu.rf_ram.memory[46][4] ;
 wire \u_cpu.rf_ram.memory[46][5] ;
 wire \u_cpu.rf_ram.memory[46][6] ;
 wire \u_cpu.rf_ram.memory[46][7] ;
 wire \u_cpu.rf_ram.memory[47][0] ;
 wire \u_cpu.rf_ram.memory[47][1] ;
 wire \u_cpu.rf_ram.memory[47][2] ;
 wire \u_cpu.rf_ram.memory[47][3] ;
 wire \u_cpu.rf_ram.memory[47][4] ;
 wire \u_cpu.rf_ram.memory[47][5] ;
 wire \u_cpu.rf_ram.memory[47][6] ;
 wire \u_cpu.rf_ram.memory[47][7] ;
 wire \u_cpu.rf_ram.memory[48][0] ;
 wire \u_cpu.rf_ram.memory[48][1] ;
 wire \u_cpu.rf_ram.memory[48][2] ;
 wire \u_cpu.rf_ram.memory[48][3] ;
 wire \u_cpu.rf_ram.memory[48][4] ;
 wire \u_cpu.rf_ram.memory[48][5] ;
 wire \u_cpu.rf_ram.memory[48][6] ;
 wire \u_cpu.rf_ram.memory[48][7] ;
 wire \u_cpu.rf_ram.memory[49][0] ;
 wire \u_cpu.rf_ram.memory[49][1] ;
 wire \u_cpu.rf_ram.memory[49][2] ;
 wire \u_cpu.rf_ram.memory[49][3] ;
 wire \u_cpu.rf_ram.memory[49][4] ;
 wire \u_cpu.rf_ram.memory[49][5] ;
 wire \u_cpu.rf_ram.memory[49][6] ;
 wire \u_cpu.rf_ram.memory[49][7] ;
 wire \u_cpu.rf_ram.memory[4][0] ;
 wire \u_cpu.rf_ram.memory[4][1] ;
 wire \u_cpu.rf_ram.memory[4][2] ;
 wire \u_cpu.rf_ram.memory[4][3] ;
 wire \u_cpu.rf_ram.memory[4][4] ;
 wire \u_cpu.rf_ram.memory[4][5] ;
 wire \u_cpu.rf_ram.memory[4][6] ;
 wire \u_cpu.rf_ram.memory[4][7] ;
 wire \u_cpu.rf_ram.memory[50][0] ;
 wire \u_cpu.rf_ram.memory[50][1] ;
 wire \u_cpu.rf_ram.memory[50][2] ;
 wire \u_cpu.rf_ram.memory[50][3] ;
 wire \u_cpu.rf_ram.memory[50][4] ;
 wire \u_cpu.rf_ram.memory[50][5] ;
 wire \u_cpu.rf_ram.memory[50][6] ;
 wire \u_cpu.rf_ram.memory[50][7] ;
 wire \u_cpu.rf_ram.memory[51][0] ;
 wire \u_cpu.rf_ram.memory[51][1] ;
 wire \u_cpu.rf_ram.memory[51][2] ;
 wire \u_cpu.rf_ram.memory[51][3] ;
 wire \u_cpu.rf_ram.memory[51][4] ;
 wire \u_cpu.rf_ram.memory[51][5] ;
 wire \u_cpu.rf_ram.memory[51][6] ;
 wire \u_cpu.rf_ram.memory[51][7] ;
 wire \u_cpu.rf_ram.memory[52][0] ;
 wire \u_cpu.rf_ram.memory[52][1] ;
 wire \u_cpu.rf_ram.memory[52][2] ;
 wire \u_cpu.rf_ram.memory[52][3] ;
 wire \u_cpu.rf_ram.memory[52][4] ;
 wire \u_cpu.rf_ram.memory[52][5] ;
 wire \u_cpu.rf_ram.memory[52][6] ;
 wire \u_cpu.rf_ram.memory[52][7] ;
 wire \u_cpu.rf_ram.memory[53][0] ;
 wire \u_cpu.rf_ram.memory[53][1] ;
 wire \u_cpu.rf_ram.memory[53][2] ;
 wire \u_cpu.rf_ram.memory[53][3] ;
 wire \u_cpu.rf_ram.memory[53][4] ;
 wire \u_cpu.rf_ram.memory[53][5] ;
 wire \u_cpu.rf_ram.memory[53][6] ;
 wire \u_cpu.rf_ram.memory[53][7] ;
 wire \u_cpu.rf_ram.memory[54][0] ;
 wire \u_cpu.rf_ram.memory[54][1] ;
 wire \u_cpu.rf_ram.memory[54][2] ;
 wire \u_cpu.rf_ram.memory[54][3] ;
 wire \u_cpu.rf_ram.memory[54][4] ;
 wire \u_cpu.rf_ram.memory[54][5] ;
 wire \u_cpu.rf_ram.memory[54][6] ;
 wire \u_cpu.rf_ram.memory[54][7] ;
 wire \u_cpu.rf_ram.memory[55][0] ;
 wire \u_cpu.rf_ram.memory[55][1] ;
 wire \u_cpu.rf_ram.memory[55][2] ;
 wire \u_cpu.rf_ram.memory[55][3] ;
 wire \u_cpu.rf_ram.memory[55][4] ;
 wire \u_cpu.rf_ram.memory[55][5] ;
 wire \u_cpu.rf_ram.memory[55][6] ;
 wire \u_cpu.rf_ram.memory[55][7] ;
 wire \u_cpu.rf_ram.memory[56][0] ;
 wire \u_cpu.rf_ram.memory[56][1] ;
 wire \u_cpu.rf_ram.memory[56][2] ;
 wire \u_cpu.rf_ram.memory[56][3] ;
 wire \u_cpu.rf_ram.memory[56][4] ;
 wire \u_cpu.rf_ram.memory[56][5] ;
 wire \u_cpu.rf_ram.memory[56][6] ;
 wire \u_cpu.rf_ram.memory[56][7] ;
 wire \u_cpu.rf_ram.memory[57][0] ;
 wire \u_cpu.rf_ram.memory[57][1] ;
 wire \u_cpu.rf_ram.memory[57][2] ;
 wire \u_cpu.rf_ram.memory[57][3] ;
 wire \u_cpu.rf_ram.memory[57][4] ;
 wire \u_cpu.rf_ram.memory[57][5] ;
 wire \u_cpu.rf_ram.memory[57][6] ;
 wire \u_cpu.rf_ram.memory[57][7] ;
 wire \u_cpu.rf_ram.memory[58][0] ;
 wire \u_cpu.rf_ram.memory[58][1] ;
 wire \u_cpu.rf_ram.memory[58][2] ;
 wire \u_cpu.rf_ram.memory[58][3] ;
 wire \u_cpu.rf_ram.memory[58][4] ;
 wire \u_cpu.rf_ram.memory[58][5] ;
 wire \u_cpu.rf_ram.memory[58][6] ;
 wire \u_cpu.rf_ram.memory[58][7] ;
 wire \u_cpu.rf_ram.memory[59][0] ;
 wire \u_cpu.rf_ram.memory[59][1] ;
 wire \u_cpu.rf_ram.memory[59][2] ;
 wire \u_cpu.rf_ram.memory[59][3] ;
 wire \u_cpu.rf_ram.memory[59][4] ;
 wire \u_cpu.rf_ram.memory[59][5] ;
 wire \u_cpu.rf_ram.memory[59][6] ;
 wire \u_cpu.rf_ram.memory[59][7] ;
 wire \u_cpu.rf_ram.memory[5][0] ;
 wire \u_cpu.rf_ram.memory[5][1] ;
 wire \u_cpu.rf_ram.memory[5][2] ;
 wire \u_cpu.rf_ram.memory[5][3] ;
 wire \u_cpu.rf_ram.memory[5][4] ;
 wire \u_cpu.rf_ram.memory[5][5] ;
 wire \u_cpu.rf_ram.memory[5][6] ;
 wire \u_cpu.rf_ram.memory[5][7] ;
 wire \u_cpu.rf_ram.memory[60][0] ;
 wire \u_cpu.rf_ram.memory[60][1] ;
 wire \u_cpu.rf_ram.memory[60][2] ;
 wire \u_cpu.rf_ram.memory[60][3] ;
 wire \u_cpu.rf_ram.memory[60][4] ;
 wire \u_cpu.rf_ram.memory[60][5] ;
 wire \u_cpu.rf_ram.memory[60][6] ;
 wire \u_cpu.rf_ram.memory[60][7] ;
 wire \u_cpu.rf_ram.memory[61][0] ;
 wire \u_cpu.rf_ram.memory[61][1] ;
 wire \u_cpu.rf_ram.memory[61][2] ;
 wire \u_cpu.rf_ram.memory[61][3] ;
 wire \u_cpu.rf_ram.memory[61][4] ;
 wire \u_cpu.rf_ram.memory[61][5] ;
 wire \u_cpu.rf_ram.memory[61][6] ;
 wire \u_cpu.rf_ram.memory[61][7] ;
 wire \u_cpu.rf_ram.memory[62][0] ;
 wire \u_cpu.rf_ram.memory[62][1] ;
 wire \u_cpu.rf_ram.memory[62][2] ;
 wire \u_cpu.rf_ram.memory[62][3] ;
 wire \u_cpu.rf_ram.memory[62][4] ;
 wire \u_cpu.rf_ram.memory[62][5] ;
 wire \u_cpu.rf_ram.memory[62][6] ;
 wire \u_cpu.rf_ram.memory[62][7] ;
 wire \u_cpu.rf_ram.memory[63][0] ;
 wire \u_cpu.rf_ram.memory[63][1] ;
 wire \u_cpu.rf_ram.memory[63][2] ;
 wire \u_cpu.rf_ram.memory[63][3] ;
 wire \u_cpu.rf_ram.memory[63][4] ;
 wire \u_cpu.rf_ram.memory[63][5] ;
 wire \u_cpu.rf_ram.memory[63][6] ;
 wire \u_cpu.rf_ram.memory[63][7] ;
 wire \u_cpu.rf_ram.memory[64][0] ;
 wire \u_cpu.rf_ram.memory[64][1] ;
 wire \u_cpu.rf_ram.memory[64][2] ;
 wire \u_cpu.rf_ram.memory[64][3] ;
 wire \u_cpu.rf_ram.memory[64][4] ;
 wire \u_cpu.rf_ram.memory[64][5] ;
 wire \u_cpu.rf_ram.memory[64][6] ;
 wire \u_cpu.rf_ram.memory[64][7] ;
 wire \u_cpu.rf_ram.memory[65][0] ;
 wire \u_cpu.rf_ram.memory[65][1] ;
 wire \u_cpu.rf_ram.memory[65][2] ;
 wire \u_cpu.rf_ram.memory[65][3] ;
 wire \u_cpu.rf_ram.memory[65][4] ;
 wire \u_cpu.rf_ram.memory[65][5] ;
 wire \u_cpu.rf_ram.memory[65][6] ;
 wire \u_cpu.rf_ram.memory[65][7] ;
 wire \u_cpu.rf_ram.memory[66][0] ;
 wire \u_cpu.rf_ram.memory[66][1] ;
 wire \u_cpu.rf_ram.memory[66][2] ;
 wire \u_cpu.rf_ram.memory[66][3] ;
 wire \u_cpu.rf_ram.memory[66][4] ;
 wire \u_cpu.rf_ram.memory[66][5] ;
 wire \u_cpu.rf_ram.memory[66][6] ;
 wire \u_cpu.rf_ram.memory[66][7] ;
 wire \u_cpu.rf_ram.memory[67][0] ;
 wire \u_cpu.rf_ram.memory[67][1] ;
 wire \u_cpu.rf_ram.memory[67][2] ;
 wire \u_cpu.rf_ram.memory[67][3] ;
 wire \u_cpu.rf_ram.memory[67][4] ;
 wire \u_cpu.rf_ram.memory[67][5] ;
 wire \u_cpu.rf_ram.memory[67][6] ;
 wire \u_cpu.rf_ram.memory[67][7] ;
 wire \u_cpu.rf_ram.memory[68][0] ;
 wire \u_cpu.rf_ram.memory[68][1] ;
 wire \u_cpu.rf_ram.memory[68][2] ;
 wire \u_cpu.rf_ram.memory[68][3] ;
 wire \u_cpu.rf_ram.memory[68][4] ;
 wire \u_cpu.rf_ram.memory[68][5] ;
 wire \u_cpu.rf_ram.memory[68][6] ;
 wire \u_cpu.rf_ram.memory[68][7] ;
 wire \u_cpu.rf_ram.memory[69][0] ;
 wire \u_cpu.rf_ram.memory[69][1] ;
 wire \u_cpu.rf_ram.memory[69][2] ;
 wire \u_cpu.rf_ram.memory[69][3] ;
 wire \u_cpu.rf_ram.memory[69][4] ;
 wire \u_cpu.rf_ram.memory[69][5] ;
 wire \u_cpu.rf_ram.memory[69][6] ;
 wire \u_cpu.rf_ram.memory[69][7] ;
 wire \u_cpu.rf_ram.memory[6][0] ;
 wire \u_cpu.rf_ram.memory[6][1] ;
 wire \u_cpu.rf_ram.memory[6][2] ;
 wire \u_cpu.rf_ram.memory[6][3] ;
 wire \u_cpu.rf_ram.memory[6][4] ;
 wire \u_cpu.rf_ram.memory[6][5] ;
 wire \u_cpu.rf_ram.memory[6][6] ;
 wire \u_cpu.rf_ram.memory[6][7] ;
 wire \u_cpu.rf_ram.memory[70][0] ;
 wire \u_cpu.rf_ram.memory[70][1] ;
 wire \u_cpu.rf_ram.memory[70][2] ;
 wire \u_cpu.rf_ram.memory[70][3] ;
 wire \u_cpu.rf_ram.memory[70][4] ;
 wire \u_cpu.rf_ram.memory[70][5] ;
 wire \u_cpu.rf_ram.memory[70][6] ;
 wire \u_cpu.rf_ram.memory[70][7] ;
 wire \u_cpu.rf_ram.memory[71][0] ;
 wire \u_cpu.rf_ram.memory[71][1] ;
 wire \u_cpu.rf_ram.memory[71][2] ;
 wire \u_cpu.rf_ram.memory[71][3] ;
 wire \u_cpu.rf_ram.memory[71][4] ;
 wire \u_cpu.rf_ram.memory[71][5] ;
 wire \u_cpu.rf_ram.memory[71][6] ;
 wire \u_cpu.rf_ram.memory[71][7] ;
 wire \u_cpu.rf_ram.memory[72][0] ;
 wire \u_cpu.rf_ram.memory[72][1] ;
 wire \u_cpu.rf_ram.memory[72][2] ;
 wire \u_cpu.rf_ram.memory[72][3] ;
 wire \u_cpu.rf_ram.memory[72][4] ;
 wire \u_cpu.rf_ram.memory[72][5] ;
 wire \u_cpu.rf_ram.memory[72][6] ;
 wire \u_cpu.rf_ram.memory[72][7] ;
 wire \u_cpu.rf_ram.memory[73][0] ;
 wire \u_cpu.rf_ram.memory[73][1] ;
 wire \u_cpu.rf_ram.memory[73][2] ;
 wire \u_cpu.rf_ram.memory[73][3] ;
 wire \u_cpu.rf_ram.memory[73][4] ;
 wire \u_cpu.rf_ram.memory[73][5] ;
 wire \u_cpu.rf_ram.memory[73][6] ;
 wire \u_cpu.rf_ram.memory[73][7] ;
 wire \u_cpu.rf_ram.memory[74][0] ;
 wire \u_cpu.rf_ram.memory[74][1] ;
 wire \u_cpu.rf_ram.memory[74][2] ;
 wire \u_cpu.rf_ram.memory[74][3] ;
 wire \u_cpu.rf_ram.memory[74][4] ;
 wire \u_cpu.rf_ram.memory[74][5] ;
 wire \u_cpu.rf_ram.memory[74][6] ;
 wire \u_cpu.rf_ram.memory[74][7] ;
 wire \u_cpu.rf_ram.memory[75][0] ;
 wire \u_cpu.rf_ram.memory[75][1] ;
 wire \u_cpu.rf_ram.memory[75][2] ;
 wire \u_cpu.rf_ram.memory[75][3] ;
 wire \u_cpu.rf_ram.memory[75][4] ;
 wire \u_cpu.rf_ram.memory[75][5] ;
 wire \u_cpu.rf_ram.memory[75][6] ;
 wire \u_cpu.rf_ram.memory[75][7] ;
 wire \u_cpu.rf_ram.memory[76][0] ;
 wire \u_cpu.rf_ram.memory[76][1] ;
 wire \u_cpu.rf_ram.memory[76][2] ;
 wire \u_cpu.rf_ram.memory[76][3] ;
 wire \u_cpu.rf_ram.memory[76][4] ;
 wire \u_cpu.rf_ram.memory[76][5] ;
 wire \u_cpu.rf_ram.memory[76][6] ;
 wire \u_cpu.rf_ram.memory[76][7] ;
 wire \u_cpu.rf_ram.memory[77][0] ;
 wire \u_cpu.rf_ram.memory[77][1] ;
 wire \u_cpu.rf_ram.memory[77][2] ;
 wire \u_cpu.rf_ram.memory[77][3] ;
 wire \u_cpu.rf_ram.memory[77][4] ;
 wire \u_cpu.rf_ram.memory[77][5] ;
 wire \u_cpu.rf_ram.memory[77][6] ;
 wire \u_cpu.rf_ram.memory[77][7] ;
 wire \u_cpu.rf_ram.memory[78][0] ;
 wire \u_cpu.rf_ram.memory[78][1] ;
 wire \u_cpu.rf_ram.memory[78][2] ;
 wire \u_cpu.rf_ram.memory[78][3] ;
 wire \u_cpu.rf_ram.memory[78][4] ;
 wire \u_cpu.rf_ram.memory[78][5] ;
 wire \u_cpu.rf_ram.memory[78][6] ;
 wire \u_cpu.rf_ram.memory[78][7] ;
 wire \u_cpu.rf_ram.memory[79][0] ;
 wire \u_cpu.rf_ram.memory[79][1] ;
 wire \u_cpu.rf_ram.memory[79][2] ;
 wire \u_cpu.rf_ram.memory[79][3] ;
 wire \u_cpu.rf_ram.memory[79][4] ;
 wire \u_cpu.rf_ram.memory[79][5] ;
 wire \u_cpu.rf_ram.memory[79][6] ;
 wire \u_cpu.rf_ram.memory[79][7] ;
 wire \u_cpu.rf_ram.memory[7][0] ;
 wire \u_cpu.rf_ram.memory[7][1] ;
 wire \u_cpu.rf_ram.memory[7][2] ;
 wire \u_cpu.rf_ram.memory[7][3] ;
 wire \u_cpu.rf_ram.memory[7][4] ;
 wire \u_cpu.rf_ram.memory[7][5] ;
 wire \u_cpu.rf_ram.memory[7][6] ;
 wire \u_cpu.rf_ram.memory[7][7] ;
 wire \u_cpu.rf_ram.memory[80][0] ;
 wire \u_cpu.rf_ram.memory[80][1] ;
 wire \u_cpu.rf_ram.memory[80][2] ;
 wire \u_cpu.rf_ram.memory[80][3] ;
 wire \u_cpu.rf_ram.memory[80][4] ;
 wire \u_cpu.rf_ram.memory[80][5] ;
 wire \u_cpu.rf_ram.memory[80][6] ;
 wire \u_cpu.rf_ram.memory[80][7] ;
 wire \u_cpu.rf_ram.memory[81][0] ;
 wire \u_cpu.rf_ram.memory[81][1] ;
 wire \u_cpu.rf_ram.memory[81][2] ;
 wire \u_cpu.rf_ram.memory[81][3] ;
 wire \u_cpu.rf_ram.memory[81][4] ;
 wire \u_cpu.rf_ram.memory[81][5] ;
 wire \u_cpu.rf_ram.memory[81][6] ;
 wire \u_cpu.rf_ram.memory[81][7] ;
 wire \u_cpu.rf_ram.memory[82][0] ;
 wire \u_cpu.rf_ram.memory[82][1] ;
 wire \u_cpu.rf_ram.memory[82][2] ;
 wire \u_cpu.rf_ram.memory[82][3] ;
 wire \u_cpu.rf_ram.memory[82][4] ;
 wire \u_cpu.rf_ram.memory[82][5] ;
 wire \u_cpu.rf_ram.memory[82][6] ;
 wire \u_cpu.rf_ram.memory[82][7] ;
 wire \u_cpu.rf_ram.memory[83][0] ;
 wire \u_cpu.rf_ram.memory[83][1] ;
 wire \u_cpu.rf_ram.memory[83][2] ;
 wire \u_cpu.rf_ram.memory[83][3] ;
 wire \u_cpu.rf_ram.memory[83][4] ;
 wire \u_cpu.rf_ram.memory[83][5] ;
 wire \u_cpu.rf_ram.memory[83][6] ;
 wire \u_cpu.rf_ram.memory[83][7] ;
 wire \u_cpu.rf_ram.memory[84][0] ;
 wire \u_cpu.rf_ram.memory[84][1] ;
 wire \u_cpu.rf_ram.memory[84][2] ;
 wire \u_cpu.rf_ram.memory[84][3] ;
 wire \u_cpu.rf_ram.memory[84][4] ;
 wire \u_cpu.rf_ram.memory[84][5] ;
 wire \u_cpu.rf_ram.memory[84][6] ;
 wire \u_cpu.rf_ram.memory[84][7] ;
 wire \u_cpu.rf_ram.memory[85][0] ;
 wire \u_cpu.rf_ram.memory[85][1] ;
 wire \u_cpu.rf_ram.memory[85][2] ;
 wire \u_cpu.rf_ram.memory[85][3] ;
 wire \u_cpu.rf_ram.memory[85][4] ;
 wire \u_cpu.rf_ram.memory[85][5] ;
 wire \u_cpu.rf_ram.memory[85][6] ;
 wire \u_cpu.rf_ram.memory[85][7] ;
 wire \u_cpu.rf_ram.memory[86][0] ;
 wire \u_cpu.rf_ram.memory[86][1] ;
 wire \u_cpu.rf_ram.memory[86][2] ;
 wire \u_cpu.rf_ram.memory[86][3] ;
 wire \u_cpu.rf_ram.memory[86][4] ;
 wire \u_cpu.rf_ram.memory[86][5] ;
 wire \u_cpu.rf_ram.memory[86][6] ;
 wire \u_cpu.rf_ram.memory[86][7] ;
 wire \u_cpu.rf_ram.memory[87][0] ;
 wire \u_cpu.rf_ram.memory[87][1] ;
 wire \u_cpu.rf_ram.memory[87][2] ;
 wire \u_cpu.rf_ram.memory[87][3] ;
 wire \u_cpu.rf_ram.memory[87][4] ;
 wire \u_cpu.rf_ram.memory[87][5] ;
 wire \u_cpu.rf_ram.memory[87][6] ;
 wire \u_cpu.rf_ram.memory[87][7] ;
 wire \u_cpu.rf_ram.memory[88][0] ;
 wire \u_cpu.rf_ram.memory[88][1] ;
 wire \u_cpu.rf_ram.memory[88][2] ;
 wire \u_cpu.rf_ram.memory[88][3] ;
 wire \u_cpu.rf_ram.memory[88][4] ;
 wire \u_cpu.rf_ram.memory[88][5] ;
 wire \u_cpu.rf_ram.memory[88][6] ;
 wire \u_cpu.rf_ram.memory[88][7] ;
 wire \u_cpu.rf_ram.memory[89][0] ;
 wire \u_cpu.rf_ram.memory[89][1] ;
 wire \u_cpu.rf_ram.memory[89][2] ;
 wire \u_cpu.rf_ram.memory[89][3] ;
 wire \u_cpu.rf_ram.memory[89][4] ;
 wire \u_cpu.rf_ram.memory[89][5] ;
 wire \u_cpu.rf_ram.memory[89][6] ;
 wire \u_cpu.rf_ram.memory[89][7] ;
 wire \u_cpu.rf_ram.memory[8][0] ;
 wire \u_cpu.rf_ram.memory[8][1] ;
 wire \u_cpu.rf_ram.memory[8][2] ;
 wire \u_cpu.rf_ram.memory[8][3] ;
 wire \u_cpu.rf_ram.memory[8][4] ;
 wire \u_cpu.rf_ram.memory[8][5] ;
 wire \u_cpu.rf_ram.memory[8][6] ;
 wire \u_cpu.rf_ram.memory[8][7] ;
 wire \u_cpu.rf_ram.memory[90][0] ;
 wire \u_cpu.rf_ram.memory[90][1] ;
 wire \u_cpu.rf_ram.memory[90][2] ;
 wire \u_cpu.rf_ram.memory[90][3] ;
 wire \u_cpu.rf_ram.memory[90][4] ;
 wire \u_cpu.rf_ram.memory[90][5] ;
 wire \u_cpu.rf_ram.memory[90][6] ;
 wire \u_cpu.rf_ram.memory[90][7] ;
 wire \u_cpu.rf_ram.memory[91][0] ;
 wire \u_cpu.rf_ram.memory[91][1] ;
 wire \u_cpu.rf_ram.memory[91][2] ;
 wire \u_cpu.rf_ram.memory[91][3] ;
 wire \u_cpu.rf_ram.memory[91][4] ;
 wire \u_cpu.rf_ram.memory[91][5] ;
 wire \u_cpu.rf_ram.memory[91][6] ;
 wire \u_cpu.rf_ram.memory[91][7] ;
 wire \u_cpu.rf_ram.memory[92][0] ;
 wire \u_cpu.rf_ram.memory[92][1] ;
 wire \u_cpu.rf_ram.memory[92][2] ;
 wire \u_cpu.rf_ram.memory[92][3] ;
 wire \u_cpu.rf_ram.memory[92][4] ;
 wire \u_cpu.rf_ram.memory[92][5] ;
 wire \u_cpu.rf_ram.memory[92][6] ;
 wire \u_cpu.rf_ram.memory[92][7] ;
 wire \u_cpu.rf_ram.memory[93][0] ;
 wire \u_cpu.rf_ram.memory[93][1] ;
 wire \u_cpu.rf_ram.memory[93][2] ;
 wire \u_cpu.rf_ram.memory[93][3] ;
 wire \u_cpu.rf_ram.memory[93][4] ;
 wire \u_cpu.rf_ram.memory[93][5] ;
 wire \u_cpu.rf_ram.memory[93][6] ;
 wire \u_cpu.rf_ram.memory[93][7] ;
 wire \u_cpu.rf_ram.memory[94][0] ;
 wire \u_cpu.rf_ram.memory[94][1] ;
 wire \u_cpu.rf_ram.memory[94][2] ;
 wire \u_cpu.rf_ram.memory[94][3] ;
 wire \u_cpu.rf_ram.memory[94][4] ;
 wire \u_cpu.rf_ram.memory[94][5] ;
 wire \u_cpu.rf_ram.memory[94][6] ;
 wire \u_cpu.rf_ram.memory[94][7] ;
 wire \u_cpu.rf_ram.memory[95][0] ;
 wire \u_cpu.rf_ram.memory[95][1] ;
 wire \u_cpu.rf_ram.memory[95][2] ;
 wire \u_cpu.rf_ram.memory[95][3] ;
 wire \u_cpu.rf_ram.memory[95][4] ;
 wire \u_cpu.rf_ram.memory[95][5] ;
 wire \u_cpu.rf_ram.memory[95][6] ;
 wire \u_cpu.rf_ram.memory[95][7] ;
 wire \u_cpu.rf_ram.memory[96][0] ;
 wire \u_cpu.rf_ram.memory[96][1] ;
 wire \u_cpu.rf_ram.memory[96][2] ;
 wire \u_cpu.rf_ram.memory[96][3] ;
 wire \u_cpu.rf_ram.memory[96][4] ;
 wire \u_cpu.rf_ram.memory[96][5] ;
 wire \u_cpu.rf_ram.memory[96][6] ;
 wire \u_cpu.rf_ram.memory[96][7] ;
 wire \u_cpu.rf_ram.memory[97][0] ;
 wire \u_cpu.rf_ram.memory[97][1] ;
 wire \u_cpu.rf_ram.memory[97][2] ;
 wire \u_cpu.rf_ram.memory[97][3] ;
 wire \u_cpu.rf_ram.memory[97][4] ;
 wire \u_cpu.rf_ram.memory[97][5] ;
 wire \u_cpu.rf_ram.memory[97][6] ;
 wire \u_cpu.rf_ram.memory[97][7] ;
 wire \u_cpu.rf_ram.memory[98][0] ;
 wire \u_cpu.rf_ram.memory[98][1] ;
 wire \u_cpu.rf_ram.memory[98][2] ;
 wire \u_cpu.rf_ram.memory[98][3] ;
 wire \u_cpu.rf_ram.memory[98][4] ;
 wire \u_cpu.rf_ram.memory[98][5] ;
 wire \u_cpu.rf_ram.memory[98][6] ;
 wire \u_cpu.rf_ram.memory[98][7] ;
 wire \u_cpu.rf_ram.memory[99][0] ;
 wire \u_cpu.rf_ram.memory[99][1] ;
 wire \u_cpu.rf_ram.memory[99][2] ;
 wire \u_cpu.rf_ram.memory[99][3] ;
 wire \u_cpu.rf_ram.memory[99][4] ;
 wire \u_cpu.rf_ram.memory[99][5] ;
 wire \u_cpu.rf_ram.memory[99][6] ;
 wire \u_cpu.rf_ram.memory[99][7] ;
 wire \u_cpu.rf_ram.memory[9][0] ;
 wire \u_cpu.rf_ram.memory[9][1] ;
 wire \u_cpu.rf_ram.memory[9][2] ;
 wire \u_cpu.rf_ram.memory[9][3] ;
 wire \u_cpu.rf_ram.memory[9][4] ;
 wire \u_cpu.rf_ram.memory[9][5] ;
 wire \u_cpu.rf_ram.memory[9][6] ;
 wire \u_cpu.rf_ram.memory[9][7] ;
 wire \u_cpu.rf_ram.rdata[0] ;
 wire \u_cpu.rf_ram.rdata[1] ;
 wire \u_cpu.rf_ram.rdata[2] ;
 wire \u_cpu.rf_ram.rdata[3] ;
 wire \u_cpu.rf_ram.rdata[4] ;
 wire \u_cpu.rf_ram.rdata[5] ;
 wire \u_cpu.rf_ram.rdata[6] ;
 wire \u_cpu.rf_ram.rdata[7] ;
 wire \u_cpu.rf_ram.regzero ;
 wire \u_cpu.rf_ram_if.genblk1.wtrig0_r ;
 wire \u_cpu.rf_ram_if.rcnt[0] ;
 wire \u_cpu.rf_ram_if.rcnt[1] ;
 wire \u_cpu.rf_ram_if.rcnt[2] ;
 wire \u_cpu.rf_ram_if.rdata0[1] ;
 wire \u_cpu.rf_ram_if.rdata0[2] ;
 wire \u_cpu.rf_ram_if.rdata0[3] ;
 wire \u_cpu.rf_ram_if.rdata0[4] ;
 wire \u_cpu.rf_ram_if.rdata0[5] ;
 wire \u_cpu.rf_ram_if.rdata0[6] ;
 wire \u_cpu.rf_ram_if.rdata0[7] ;
 wire \u_cpu.rf_ram_if.rdata1[0] ;
 wire \u_cpu.rf_ram_if.rdata1[1] ;
 wire \u_cpu.rf_ram_if.rdata1[2] ;
 wire \u_cpu.rf_ram_if.rdata1[3] ;
 wire \u_cpu.rf_ram_if.rdata1[4] ;
 wire \u_cpu.rf_ram_if.rdata1[5] ;
 wire \u_cpu.rf_ram_if.rdata1[6] ;
 wire \u_cpu.rf_ram_if.rgnt ;
 wire \u_cpu.rf_ram_if.rreq_r ;
 wire \u_cpu.rf_ram_if.rtrig0 ;
 wire \u_cpu.rf_ram_if.rtrig1 ;
 wire \u_cpu.rf_ram_if.wdata0_r[0] ;
 wire \u_cpu.rf_ram_if.wdata0_r[1] ;
 wire \u_cpu.rf_ram_if.wdata0_r[2] ;
 wire \u_cpu.rf_ram_if.wdata0_r[3] ;
 wire \u_cpu.rf_ram_if.wdata0_r[4] ;
 wire \u_cpu.rf_ram_if.wdata0_r[5] ;
 wire \u_cpu.rf_ram_if.wdata0_r[6] ;
 wire \u_cpu.rf_ram_if.wdata1_r[0] ;
 wire \u_cpu.rf_ram_if.wdata1_r[1] ;
 wire \u_cpu.rf_ram_if.wdata1_r[2] ;
 wire \u_cpu.rf_ram_if.wdata1_r[3] ;
 wire \u_cpu.rf_ram_if.wdata1_r[4] ;
 wire \u_cpu.rf_ram_if.wdata1_r[5] ;
 wire \u_cpu.rf_ram_if.wdata1_r[6] ;
 wire \u_cpu.rf_ram_if.wdata1_r[7] ;
 wire \u_cpu.rf_ram_if.wen0_r ;
 wire \u_cpu.rf_ram_if.wen1_r ;
 wire \u_cpu.rf_ram_if.wtrig0 ;
 wire \u_scanchain_local.data_out ;
 wire \u_scanchain_local.module_data_in[34] ;
 wire \u_scanchain_local.module_data_in[35] ;
 wire \u_scanchain_local.module_data_in[36] ;
 wire \u_scanchain_local.module_data_in[37] ;
 wire \u_scanchain_local.module_data_in[38] ;
 wire \u_scanchain_local.module_data_in[39] ;
 wire \u_scanchain_local.module_data_in[40] ;
 wire \u_scanchain_local.module_data_in[41] ;
 wire \u_scanchain_local.module_data_in[42] ;
 wire \u_scanchain_local.module_data_in[43] ;
 wire \u_scanchain_local.module_data_in[44] ;
 wire \u_scanchain_local.module_data_in[45] ;
 wire \u_scanchain_local.module_data_in[46] ;
 wire \u_scanchain_local.module_data_in[47] ;
 wire \u_scanchain_local.module_data_in[48] ;
 wire \u_scanchain_local.module_data_in[49] ;
 wire \u_scanchain_local.module_data_in[50] ;
 wire \u_scanchain_local.module_data_in[51] ;
 wire \u_scanchain_local.module_data_in[52] ;
 wire \u_scanchain_local.module_data_in[53] ;
 wire \u_scanchain_local.module_data_in[54] ;
 wire \u_scanchain_local.module_data_in[55] ;
 wire \u_scanchain_local.module_data_in[56] ;
 wire \u_scanchain_local.module_data_in[57] ;
 wire \u_scanchain_local.module_data_in[58] ;
 wire \u_scanchain_local.module_data_in[59] ;
 wire \u_scanchain_local.module_data_in[60] ;
 wire \u_scanchain_local.module_data_in[61] ;
 wire \u_scanchain_local.module_data_in[62] ;
 wire \u_scanchain_local.module_data_in[63] ;
 wire \u_scanchain_local.module_data_in[64] ;
 wire \u_scanchain_local.module_data_in[65] ;
 wire \u_scanchain_local.module_data_in[66] ;
 wire \u_scanchain_local.module_data_in[67] ;
 wire \u_scanchain_local.module_data_in[68] ;
 wire \u_scanchain_local.module_data_in[69] ;

 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _04848_ (.I(\u_cpu.rf_ram_if.rcnt[0] ),
    .ZN(_01436_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _04849_ (.A1(_01436_),
    .A2(\u_cpu.rf_ram_if.rcnt[2] ),
    .A3(\u_cpu.rf_ram_if.rcnt[1] ),
    .Z(_01437_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _04850_ (.I(_01437_),
    .Z(_01438_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _04851_ (.I(_01438_),
    .ZN(\u_cpu.rf_ram_if.rtrig0 ));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _04852_ (.I(\u_cpu.cpu.csr_imm ),
    .ZN(_01439_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _04853_ (.I(\u_cpu.cpu.immdec.imm24_20[0] ),
    .ZN(_01440_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _04854_ (.I(\u_cpu.cpu.decode.co_mem_word ),
    .Z(_01441_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _04855_ (.I(\u_cpu.cpu.csr_d_sel ),
    .Z(_01442_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _04856_ (.A1(_01441_),
    .A2(\u_cpu.cpu.bne_or_bge ),
    .A3(_01442_),
    .Z(_01443_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _04857_ (.I(\u_cpu.cpu.decode.opcode[2] ),
    .Z(_01444_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _04858_ (.I(\u_cpu.cpu.branch_op ),
    .Z(_01445_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _04859_ (.A1(_01444_),
    .A2(_01445_),
    .Z(_01446_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _04860_ (.A1(_01443_),
    .A2(_01446_),
    .ZN(_01447_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _04861_ (.I(\u_cpu.cpu.decode.op21 ),
    .ZN(_01448_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _04862_ (.A1(_01448_),
    .A2(\u_cpu.cpu.decode.op26 ),
    .B(\u_cpu.cpu.decode.co_ebreak ),
    .ZN(_01449_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _04863_ (.A1(_01441_),
    .A2(\u_cpu.cpu.bne_or_bge ),
    .A3(_01442_),
    .ZN(_01450_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _04864_ (.A1(_01450_),
    .A2(_01446_),
    .B(\u_cpu.cpu.genblk3.csr.o_new_irq ),
    .C(\u_cpu.cpu.state.genblk1.misalign_trap_sync_r ),
    .ZN(_01451_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _04865_ (.A1(_01447_),
    .A2(_01449_),
    .B(_01451_),
    .ZN(_01452_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _04866_ (.A1(_01440_),
    .A2(_01452_),
    .ZN(_01453_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _04867_ (.I(\u_cpu.cpu.decode.op26 ),
    .ZN(_01454_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _04868_ (.A1(\u_cpu.cpu.decode.op21 ),
    .A2(_01454_),
    .ZN(_01455_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _04869_ (.A1(_01447_),
    .A2(_01449_),
    .Z(_01456_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _04870_ (.A1(_01444_),
    .A2(_01445_),
    .ZN(_01457_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _04871_ (.I(\u_cpu.cpu.genblk3.csr.o_new_irq ),
    .ZN(_01458_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _04872_ (.A1(\u_cpu.cpu.decode.op21 ),
    .A2(_01443_),
    .A3(_01457_),
    .B(_01458_),
    .ZN(_01459_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _04873_ (.A1(\u_cpu.cpu.state.genblk1.misalign_trap_sync_r ),
    .A2(_01459_),
    .ZN(_01460_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _04874_ (.A1(_01455_),
    .A2(_01456_),
    .B(\u_cpu.rf_ram_if.rtrig0 ),
    .C(_01460_),
    .ZN(_01461_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _04875_ (.A1(_01453_),
    .A2(_01461_),
    .ZN(_01462_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _04876_ (.A1(_01439_),
    .A2(_01438_),
    .B(_01462_),
    .ZN(_01463_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _04877_ (.I(_01463_),
    .Z(_01464_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _04878_ (.I(_01464_),
    .Z(_01465_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _04879_ (.A1(\u_cpu.rf_ram_if.rtrig0 ),
    .A2(_01452_),
    .Z(_01466_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _04880_ (.I(_01438_),
    .Z(_01467_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _04881_ (.A1(\u_cpu.cpu.immdec.imm19_12_20[8] ),
    .A2(_01467_),
    .ZN(_01468_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _04882_ (.A1(_01438_),
    .A2(_01452_),
    .ZN(_01469_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _04883_ (.A1(\u_cpu.cpu.immdec.imm24_20[4] ),
    .A2(_01469_),
    .ZN(_01470_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _04884_ (.A1(_01468_),
    .A2(_01470_),
    .ZN(_01471_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _04885_ (.A1(_01466_),
    .A2(_01471_),
    .ZN(_01472_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _04886_ (.I(_01472_),
    .Z(_01473_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _04887_ (.A1(\u_cpu.cpu.immdec.imm19_12_20[5] ),
    .A2(\u_cpu.rf_ram_if.rtrig0 ),
    .Z(_01474_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _04888_ (.I(\u_cpu.cpu.immdec.imm24_20[1] ),
    .ZN(_01475_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _04889_ (.A1(\u_cpu.cpu.decode.op26 ),
    .A2(\u_cpu.cpu.decode.co_ebreak ),
    .ZN(_01476_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _04890_ (.A1(_01448_),
    .A2(_01443_),
    .A3(_01457_),
    .ZN(_01477_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _04891_ (.A1(_01438_),
    .A2(_01477_),
    .ZN(_01478_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _04892_ (.A1(_01475_),
    .A2(_01452_),
    .B1(_01476_),
    .B2(_01447_),
    .C(_01478_),
    .ZN(_01479_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _04893_ (.A1(_01474_),
    .A2(_01479_),
    .ZN(_01480_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _04894_ (.I(_01480_),
    .Z(_01481_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _04895_ (.I(_01481_),
    .Z(_01482_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _04896_ (.A1(\u_cpu.cpu.immdec.imm19_12_20[6] ),
    .A2(_01438_),
    .ZN(_01483_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _04897_ (.A1(\u_cpu.cpu.immdec.imm24_20[2] ),
    .A2(_01469_),
    .ZN(_01484_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _04898_ (.A1(_01483_),
    .A2(_01484_),
    .Z(_01485_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _04899_ (.I(_01485_),
    .Z(_01486_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _04900_ (.A1(\u_cpu.cpu.immdec.imm19_12_20[7] ),
    .A2(_01438_),
    .ZN(_01487_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _04901_ (.A1(\u_cpu.cpu.immdec.imm24_20[3] ),
    .A2(_01469_),
    .ZN(_01488_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _04902_ (.A1(_01487_),
    .A2(_01488_),
    .Z(_01489_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _04903_ (.I(_01489_),
    .Z(_01490_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _04904_ (.A1(_01473_),
    .A2(_01482_),
    .A3(_01486_),
    .A4(_01490_),
    .ZN(_01491_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _04905_ (.A1(_01465_),
    .A2(_01491_),
    .ZN(_00025_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _04906_ (.I(_01467_),
    .ZN(\u_cpu.rf_ram_if.wtrig0 ));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _04907_ (.A1(_01487_),
    .A2(_01488_),
    .ZN(_01492_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _04908_ (.I(_01464_),
    .Z(_01493_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _04909_ (.I(\u_cpu.raddr[0] ),
    .Z(_01494_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _04910_ (.I(_01494_),
    .Z(_01495_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _04911_ (.I(_01495_),
    .Z(_01496_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _04912_ (.I(_01496_),
    .Z(_01497_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _04913_ (.I(\u_cpu.raddr[1] ),
    .Z(_01498_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _04914_ (.I(_01498_),
    .Z(_01499_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _04915_ (.I(_01499_),
    .Z(_01500_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _04916_ (.I(_01500_),
    .Z(_01501_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _04917_ (.I0(\u_cpu.rf_ram.memory[28][0] ),
    .I1(\u_cpu.rf_ram.memory[29][0] ),
    .I2(\u_cpu.rf_ram.memory[30][0] ),
    .I3(\u_cpu.rf_ram.memory[31][0] ),
    .S0(_01497_),
    .S1(_01501_),
    .Z(_01502_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _04918_ (.A1(_01493_),
    .A2(_01502_),
    .ZN(_01503_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _04919_ (.A1(\u_cpu.cpu.csr_imm ),
    .A2(\u_cpu.rf_ram_if.rtrig0 ),
    .B1(_01453_),
    .B2(_01461_),
    .ZN(_01504_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _04920_ (.I(_01504_),
    .Z(_01505_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _04921_ (.I(_01505_),
    .Z(_01506_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _04922_ (.I(_01494_),
    .Z(_01507_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _04923_ (.I(_01507_),
    .Z(_01508_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _04924_ (.I(_01499_),
    .Z(_01509_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _04925_ (.I0(\u_cpu.rf_ram.memory[24][0] ),
    .I1(\u_cpu.rf_ram.memory[25][0] ),
    .I2(\u_cpu.rf_ram.memory[26][0] ),
    .I3(\u_cpu.rf_ram.memory[27][0] ),
    .S0(_01508_),
    .S1(_01509_),
    .Z(_01510_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _04926_ (.A1(_01506_),
    .A2(_01510_),
    .B(_01481_),
    .ZN(_01511_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _04927_ (.I(_01463_),
    .Z(_01512_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _04928_ (.I(_01512_),
    .Z(_01513_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _04929_ (.I0(\u_cpu.rf_ram.memory[20][0] ),
    .I1(\u_cpu.rf_ram.memory[21][0] ),
    .I2(\u_cpu.rf_ram.memory[22][0] ),
    .I3(\u_cpu.rf_ram.memory[23][0] ),
    .S0(_01497_),
    .S1(_01501_),
    .Z(_01514_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _04930_ (.A1(_01513_),
    .A2(_01514_),
    .ZN(_01515_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _04931_ (.I0(\u_cpu.rf_ram.memory[16][0] ),
    .I1(\u_cpu.rf_ram.memory[17][0] ),
    .I2(\u_cpu.rf_ram.memory[18][0] ),
    .I3(\u_cpu.rf_ram.memory[19][0] ),
    .S0(_01508_),
    .S1(_01509_),
    .Z(_01516_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _04932_ (.A1(_01474_),
    .A2(_01479_),
    .Z(_01517_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _04933_ (.I(_01517_),
    .Z(_01518_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _04934_ (.I(_01518_),
    .Z(_01519_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _04935_ (.A1(_01506_),
    .A2(_01516_),
    .B(_01519_),
    .ZN(_01520_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _04936_ (.A1(_01503_),
    .A2(_01511_),
    .B1(_01515_),
    .B2(_01520_),
    .C(_01486_),
    .ZN(_01521_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _04937_ (.I(_01495_),
    .Z(_01522_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _04938_ (.I(_01522_),
    .Z(_01523_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _04939_ (.I(_01499_),
    .Z(_01524_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _04940_ (.I(_01524_),
    .Z(_01525_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _04941_ (.I0(\u_cpu.rf_ram.memory[4][0] ),
    .I1(\u_cpu.rf_ram.memory[5][0] ),
    .I2(\u_cpu.rf_ram.memory[6][0] ),
    .I3(\u_cpu.rf_ram.memory[7][0] ),
    .S0(_01523_),
    .S1(_01525_),
    .Z(_01526_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _04942_ (.A1(_01493_),
    .A2(_01526_),
    .ZN(_01527_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _04943_ (.I(_01505_),
    .Z(_01528_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _04944_ (.I(_01494_),
    .Z(_01529_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _04945_ (.I(_01529_),
    .Z(_01530_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _04946_ (.I(_01498_),
    .Z(_01531_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _04947_ (.I(_01531_),
    .Z(_01532_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _04948_ (.I0(\u_cpu.rf_ram.memory[0][0] ),
    .I1(\u_cpu.rf_ram.memory[1][0] ),
    .I2(\u_cpu.rf_ram.memory[2][0] ),
    .I3(\u_cpu.rf_ram.memory[3][0] ),
    .S0(_01530_),
    .S1(_01532_),
    .Z(_01533_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _04949_ (.I(_01519_),
    .Z(_01534_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _04950_ (.A1(_01528_),
    .A2(_01533_),
    .B(_01534_),
    .ZN(_01535_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _04951_ (.I0(\u_cpu.rf_ram.memory[8][0] ),
    .I1(\u_cpu.rf_ram.memory[9][0] ),
    .I2(\u_cpu.rf_ram.memory[10][0] ),
    .I3(\u_cpu.rf_ram.memory[11][0] ),
    .S0(_01523_),
    .S1(_01525_),
    .Z(_01536_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _04952_ (.A1(_01528_),
    .A2(_01536_),
    .ZN(_01537_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _04953_ (.I0(\u_cpu.rf_ram.memory[12][0] ),
    .I1(\u_cpu.rf_ram.memory[13][0] ),
    .I2(\u_cpu.rf_ram.memory[14][0] ),
    .I3(\u_cpu.rf_ram.memory[15][0] ),
    .S0(_01530_),
    .S1(_01532_),
    .Z(_01538_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _04954_ (.A1(_01513_),
    .A2(_01538_),
    .B(_01482_),
    .ZN(_01539_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _04955_ (.A1(_01483_),
    .A2(_01484_),
    .ZN(_01540_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _04956_ (.I(_01540_),
    .Z(_01541_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _04957_ (.A1(_01527_),
    .A2(_01535_),
    .B1(_01537_),
    .B2(_01539_),
    .C(_01541_),
    .ZN(_01542_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _04958_ (.I(_01463_),
    .Z(_01543_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _04959_ (.I(_01495_),
    .Z(_01544_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _04960_ (.I(_01499_),
    .Z(_01545_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _04961_ (.I0(\u_cpu.rf_ram.memory[36][0] ),
    .I1(\u_cpu.rf_ram.memory[37][0] ),
    .I2(\u_cpu.rf_ram.memory[38][0] ),
    .I3(\u_cpu.rf_ram.memory[39][0] ),
    .S0(_01544_),
    .S1(_01545_),
    .Z(_01546_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _04962_ (.A1(_01543_),
    .A2(_01546_),
    .ZN(_01547_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _04963_ (.I(_01504_),
    .Z(_01548_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _04964_ (.I0(\u_cpu.rf_ram.memory[32][0] ),
    .I1(\u_cpu.rf_ram.memory[33][0] ),
    .I2(\u_cpu.rf_ram.memory[34][0] ),
    .I3(\u_cpu.rf_ram.memory[35][0] ),
    .S0(_01495_),
    .S1(_01499_),
    .Z(_01549_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _04965_ (.A1(_01548_),
    .A2(_01549_),
    .B(_01518_),
    .ZN(_01550_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _04966_ (.I(_01495_),
    .Z(_01551_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _04967_ (.I0(\u_cpu.rf_ram.memory[40][0] ),
    .I1(\u_cpu.rf_ram.memory[41][0] ),
    .I2(\u_cpu.rf_ram.memory[42][0] ),
    .I3(\u_cpu.rf_ram.memory[43][0] ),
    .S0(_01551_),
    .S1(_01524_),
    .Z(_01552_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _04968_ (.A1(_01505_),
    .A2(_01552_),
    .ZN(_01553_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _04969_ (.I(_01463_),
    .Z(_01554_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _04970_ (.I(_01494_),
    .Z(_01555_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _04971_ (.I(_01498_),
    .Z(_01556_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _04972_ (.I0(\u_cpu.rf_ram.memory[44][0] ),
    .I1(\u_cpu.rf_ram.memory[45][0] ),
    .I2(\u_cpu.rf_ram.memory[46][0] ),
    .I3(\u_cpu.rf_ram.memory[47][0] ),
    .S0(_01555_),
    .S1(_01556_),
    .Z(_01557_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _04973_ (.I(_01480_),
    .Z(_01558_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _04974_ (.A1(_01554_),
    .A2(_01557_),
    .B(_01558_),
    .ZN(_01559_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _04975_ (.I(_01540_),
    .Z(_01560_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _04976_ (.A1(_01547_),
    .A2(_01550_),
    .B1(_01553_),
    .B2(_01559_),
    .C(_01560_),
    .ZN(_01561_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _04977_ (.I(_01495_),
    .Z(_01562_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _04978_ (.I(_01499_),
    .Z(_01563_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _04979_ (.I0(\u_cpu.rf_ram.memory[60][0] ),
    .I1(\u_cpu.rf_ram.memory[61][0] ),
    .I2(\u_cpu.rf_ram.memory[62][0] ),
    .I3(\u_cpu.rf_ram.memory[63][0] ),
    .S0(_01562_),
    .S1(_01563_),
    .Z(_01564_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _04980_ (.A1(_01464_),
    .A2(_01564_),
    .ZN(_01565_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _04981_ (.I(_01504_),
    .Z(_01566_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _04982_ (.I(_01494_),
    .Z(_01567_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _04983_ (.I(_01498_),
    .Z(_01568_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _04984_ (.I0(\u_cpu.rf_ram.memory[56][0] ),
    .I1(\u_cpu.rf_ram.memory[57][0] ),
    .I2(\u_cpu.rf_ram.memory[58][0] ),
    .I3(\u_cpu.rf_ram.memory[59][0] ),
    .S0(_01567_),
    .S1(_01568_),
    .Z(_01569_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _04985_ (.A1(_01566_),
    .A2(_01569_),
    .B(_01480_),
    .ZN(_01570_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _04986_ (.I(_01463_),
    .Z(_01571_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _04987_ (.I(_01495_),
    .Z(_01572_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _04988_ (.I(_01499_),
    .Z(_01573_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _04989_ (.I0(\u_cpu.rf_ram.memory[52][0] ),
    .I1(\u_cpu.rf_ram.memory[53][0] ),
    .I2(\u_cpu.rf_ram.memory[54][0] ),
    .I3(\u_cpu.rf_ram.memory[55][0] ),
    .S0(_01572_),
    .S1(_01573_),
    .Z(_01574_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _04990_ (.A1(_01571_),
    .A2(_01574_),
    .ZN(_01575_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _04991_ (.I(_01495_),
    .Z(_01576_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _04992_ (.I(_01498_),
    .Z(_01577_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _04993_ (.I0(\u_cpu.rf_ram.memory[48][0] ),
    .I1(\u_cpu.rf_ram.memory[49][0] ),
    .I2(\u_cpu.rf_ram.memory[50][0] ),
    .I3(\u_cpu.rf_ram.memory[51][0] ),
    .S0(_01576_),
    .S1(_01577_),
    .Z(_01578_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _04994_ (.I(_01518_),
    .Z(_01579_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _04995_ (.A1(_01505_),
    .A2(_01578_),
    .B(_01579_),
    .ZN(_01580_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _04996_ (.I(_01485_),
    .Z(_01581_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _04997_ (.A1(_01565_),
    .A2(_01570_),
    .B1(_01575_),
    .B2(_01580_),
    .C(_01581_),
    .ZN(_01582_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _04998_ (.A1(_01490_),
    .A2(_01561_),
    .A3(_01582_),
    .Z(_01583_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _04999_ (.A1(_01492_),
    .A2(_01521_),
    .A3(_01542_),
    .B(_01583_),
    .ZN(_01584_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05000_ (.I0(\u_cpu.rf_ram.memory[100][0] ),
    .I1(\u_cpu.rf_ram.memory[101][0] ),
    .I2(\u_cpu.rf_ram.memory[102][0] ),
    .I3(\u_cpu.rf_ram.memory[103][0] ),
    .S0(_01572_),
    .S1(_01573_),
    .Z(_01585_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05001_ (.A1(_01571_),
    .A2(_01585_),
    .ZN(_01586_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05002_ (.I0(\u_cpu.rf_ram.memory[96][0] ),
    .I1(\u_cpu.rf_ram.memory[97][0] ),
    .I2(\u_cpu.rf_ram.memory[98][0] ),
    .I3(\u_cpu.rf_ram.memory[99][0] ),
    .S0(_01567_),
    .S1(_01568_),
    .Z(_01587_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05003_ (.A1(_01548_),
    .A2(_01587_),
    .B(_01579_),
    .ZN(_01588_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05004_ (.I0(\u_cpu.rf_ram.memory[108][0] ),
    .I1(\u_cpu.rf_ram.memory[109][0] ),
    .I2(\u_cpu.rf_ram.memory[110][0] ),
    .I3(\u_cpu.rf_ram.memory[111][0] ),
    .S0(_01551_),
    .S1(_01524_),
    .Z(_01589_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05005_ (.A1(_01512_),
    .A2(_01589_),
    .ZN(_01590_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05006_ (.I0(\u_cpu.rf_ram.memory[104][0] ),
    .I1(\u_cpu.rf_ram.memory[105][0] ),
    .I2(\u_cpu.rf_ram.memory[106][0] ),
    .I3(\u_cpu.rf_ram.memory[107][0] ),
    .S0(_01555_),
    .S1(_01531_),
    .Z(_01591_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05007_ (.A1(_01566_),
    .A2(_01591_),
    .B(_01558_),
    .ZN(_01592_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _05008_ (.A1(_01586_),
    .A2(_01588_),
    .B1(_01590_),
    .B2(_01592_),
    .C(_01560_),
    .ZN(_01593_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05009_ (.I(_01499_),
    .Z(_01594_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05010_ (.I0(\u_cpu.rf_ram.memory[124][0] ),
    .I1(\u_cpu.rf_ram.memory[125][0] ),
    .I2(\u_cpu.rf_ram.memory[126][0] ),
    .I3(\u_cpu.rf_ram.memory[127][0] ),
    .S0(_01496_),
    .S1(_01594_),
    .Z(_01595_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05011_ (.A1(_01543_),
    .A2(_01595_),
    .ZN(_01596_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05012_ (.I(_01504_),
    .Z(_01597_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05013_ (.I(_01495_),
    .Z(_01598_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05014_ (.I0(\u_cpu.rf_ram.memory[120][0] ),
    .I1(\u_cpu.rf_ram.memory[121][0] ),
    .I2(\u_cpu.rf_ram.memory[122][0] ),
    .I3(\u_cpu.rf_ram.memory[123][0] ),
    .S0(_01598_),
    .S1(_01556_),
    .Z(_01599_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05015_ (.I(_01480_),
    .Z(_01600_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05016_ (.A1(_01597_),
    .A2(_01599_),
    .B(_01600_),
    .ZN(_01601_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05017_ (.I(_01504_),
    .Z(_01602_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05018_ (.I0(\u_cpu.rf_ram.memory[112][0] ),
    .I1(\u_cpu.rf_ram.memory[113][0] ),
    .I2(\u_cpu.rf_ram.memory[114][0] ),
    .I3(\u_cpu.rf_ram.memory[115][0] ),
    .S0(_01544_),
    .S1(_01545_),
    .Z(_01603_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05019_ (.A1(_01602_),
    .A2(_01603_),
    .ZN(_01604_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05020_ (.I(_01498_),
    .Z(_01605_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05021_ (.I0(\u_cpu.rf_ram.memory[116][0] ),
    .I1(\u_cpu.rf_ram.memory[117][0] ),
    .I2(\u_cpu.rf_ram.memory[118][0] ),
    .I3(\u_cpu.rf_ram.memory[119][0] ),
    .S0(_01576_),
    .S1(_01605_),
    .Z(_01606_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05022_ (.I(_01518_),
    .Z(_01607_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05023_ (.A1(_01554_),
    .A2(_01606_),
    .B(_01607_),
    .ZN(_01608_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _05024_ (.A1(_01596_),
    .A2(_01601_),
    .B1(_01604_),
    .B2(_01608_),
    .C(_01581_),
    .ZN(_01609_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _05025_ (.A1(_01490_),
    .A2(_01593_),
    .A3(_01609_),
    .ZN(_01610_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05026_ (.I0(\u_cpu.rf_ram.memory[92][0] ),
    .I1(\u_cpu.rf_ram.memory[93][0] ),
    .I2(\u_cpu.rf_ram.memory[94][0] ),
    .I3(\u_cpu.rf_ram.memory[95][0] ),
    .S0(_01562_),
    .S1(_01563_),
    .Z(_01611_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05027_ (.A1(_01464_),
    .A2(_01611_),
    .ZN(_01612_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05028_ (.I0(\u_cpu.rf_ram.memory[88][0] ),
    .I1(\u_cpu.rf_ram.memory[89][0] ),
    .I2(\u_cpu.rf_ram.memory[90][0] ),
    .I3(\u_cpu.rf_ram.memory[91][0] ),
    .S0(_01598_),
    .S1(_01577_),
    .Z(_01613_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05029_ (.A1(_01597_),
    .A2(_01613_),
    .B(_01600_),
    .ZN(_01614_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05030_ (.I0(\u_cpu.rf_ram.memory[80][0] ),
    .I1(\u_cpu.rf_ram.memory[81][0] ),
    .I2(\u_cpu.rf_ram.memory[82][0] ),
    .I3(\u_cpu.rf_ram.memory[83][0] ),
    .S0(_01496_),
    .S1(_01594_),
    .Z(_01615_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05031_ (.A1(_01602_),
    .A2(_01615_),
    .ZN(_01616_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05032_ (.I(_01463_),
    .Z(_01617_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05033_ (.I0(\u_cpu.rf_ram.memory[84][0] ),
    .I1(\u_cpu.rf_ram.memory[85][0] ),
    .I2(\u_cpu.rf_ram.memory[86][0] ),
    .I3(\u_cpu.rf_ram.memory[87][0] ),
    .S0(_01507_),
    .S1(_01605_),
    .Z(_01618_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05034_ (.A1(_01617_),
    .A2(_01618_),
    .B(_01607_),
    .ZN(_01619_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _05035_ (.A1(_01612_),
    .A2(_01614_),
    .B1(_01616_),
    .B2(_01619_),
    .C(_01486_),
    .ZN(_01620_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05036_ (.I(_01504_),
    .Z(_01621_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05037_ (.I(_01499_),
    .Z(_01622_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05038_ (.I0(\u_cpu.rf_ram.memory[64][0] ),
    .I1(\u_cpu.rf_ram.memory[65][0] ),
    .I2(\u_cpu.rf_ram.memory[66][0] ),
    .I3(\u_cpu.rf_ram.memory[67][0] ),
    .S0(_01522_),
    .S1(_01622_),
    .Z(_01623_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05039_ (.A1(_01621_),
    .A2(_01623_),
    .ZN(_01624_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05040_ (.I0(\u_cpu.rf_ram.memory[68][0] ),
    .I1(\u_cpu.rf_ram.memory[69][0] ),
    .I2(\u_cpu.rf_ram.memory[70][0] ),
    .I3(\u_cpu.rf_ram.memory[71][0] ),
    .S0(_01529_),
    .S1(_01500_),
    .Z(_01625_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05041_ (.A1(_01617_),
    .A2(_01625_),
    .B(_01519_),
    .ZN(_01626_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05042_ (.I0(\u_cpu.rf_ram.memory[72][0] ),
    .I1(\u_cpu.rf_ram.memory[73][0] ),
    .I2(\u_cpu.rf_ram.memory[74][0] ),
    .I3(\u_cpu.rf_ram.memory[75][0] ),
    .S0(_01522_),
    .S1(_01622_),
    .Z(_01627_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05043_ (.A1(_01621_),
    .A2(_01627_),
    .ZN(_01628_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05044_ (.I0(\u_cpu.rf_ram.memory[76][0] ),
    .I1(\u_cpu.rf_ram.memory[77][0] ),
    .I2(\u_cpu.rf_ram.memory[78][0] ),
    .I3(\u_cpu.rf_ram.memory[79][0] ),
    .S0(_01529_),
    .S1(_01500_),
    .Z(_01629_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05045_ (.A1(_01512_),
    .A2(_01629_),
    .B(_01481_),
    .ZN(_01630_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _05046_ (.A1(_01624_),
    .A2(_01626_),
    .B1(_01628_),
    .B2(_01630_),
    .C(_01541_),
    .ZN(_01631_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _05047_ (.A1(_01492_),
    .A2(_01620_),
    .A3(_01631_),
    .ZN(_01632_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05048_ (.A1(_01610_),
    .A2(_01632_),
    .B(_01471_),
    .ZN(_01633_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05049_ (.I(_01522_),
    .Z(_01634_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05050_ (.I(_01622_),
    .Z(_01635_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05051_ (.I0(\u_cpu.rf_ram.memory[136][0] ),
    .I1(\u_cpu.rf_ram.memory[137][0] ),
    .I2(\u_cpu.rf_ram.memory[138][0] ),
    .I3(\u_cpu.rf_ram.memory[139][0] ),
    .S0(_01634_),
    .S1(_01635_),
    .Z(_01636_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05052_ (.A1(_01465_),
    .A2(_01636_),
    .ZN(_01637_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05053_ (.I(_01621_),
    .Z(_01638_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05054_ (.I0(\u_cpu.rf_ram.memory[140][0] ),
    .I1(\u_cpu.rf_ram.memory[141][0] ),
    .I2(\u_cpu.rf_ram.memory[142][0] ),
    .I3(\u_cpu.rf_ram.memory[143][0] ),
    .S0(_01634_),
    .S1(_01635_),
    .Z(_01639_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05055_ (.A1(_01638_),
    .A2(_01639_),
    .B(_01534_),
    .ZN(_01640_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05056_ (.I(_01522_),
    .Z(_01641_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05057_ (.I(_01622_),
    .Z(_01642_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05058_ (.I0(\u_cpu.rf_ram.memory[128][0] ),
    .I1(\u_cpu.rf_ram.memory[129][0] ),
    .I2(\u_cpu.rf_ram.memory[130][0] ),
    .I3(\u_cpu.rf_ram.memory[131][0] ),
    .S0(_01641_),
    .S1(_01642_),
    .Z(_01643_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05059_ (.A1(_01465_),
    .A2(_01643_),
    .ZN(_01644_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05060_ (.I0(\u_cpu.rf_ram.memory[132][0] ),
    .I1(\u_cpu.rf_ram.memory[133][0] ),
    .I2(\u_cpu.rf_ram.memory[134][0] ),
    .I3(\u_cpu.rf_ram.memory[135][0] ),
    .S0(_01641_),
    .S1(_01642_),
    .Z(_01645_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05061_ (.A1(_01638_),
    .A2(_01645_),
    .B(_01482_),
    .ZN(_01646_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _05062_ (.A1(_01637_),
    .A2(_01640_),
    .B1(_01644_),
    .B2(_01646_),
    .C(_01466_),
    .ZN(_01647_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05063_ (.A1(_01633_),
    .A2(_01647_),
    .ZN(_01648_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05064_ (.A1(_01473_),
    .A2(_01584_),
    .B(_01648_),
    .ZN(_00000_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05065_ (.I0(\u_cpu.rf_ram.memory[28][1] ),
    .I1(\u_cpu.rf_ram.memory[29][1] ),
    .I2(\u_cpu.rf_ram.memory[30][1] ),
    .I3(\u_cpu.rf_ram.memory[31][1] ),
    .S0(_01497_),
    .S1(_01501_),
    .Z(_01649_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05066_ (.A1(_01493_),
    .A2(_01649_),
    .ZN(_01650_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05067_ (.I0(\u_cpu.rf_ram.memory[24][1] ),
    .I1(\u_cpu.rf_ram.memory[25][1] ),
    .I2(\u_cpu.rf_ram.memory[26][1] ),
    .I3(\u_cpu.rf_ram.memory[27][1] ),
    .S0(_01508_),
    .S1(_01509_),
    .Z(_01651_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05068_ (.A1(_01506_),
    .A2(_01651_),
    .B(_01481_),
    .ZN(_01652_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05069_ (.I0(\u_cpu.rf_ram.memory[20][1] ),
    .I1(\u_cpu.rf_ram.memory[21][1] ),
    .I2(\u_cpu.rf_ram.memory[22][1] ),
    .I3(\u_cpu.rf_ram.memory[23][1] ),
    .S0(_01497_),
    .S1(_01501_),
    .Z(_01653_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05070_ (.A1(_01513_),
    .A2(_01653_),
    .ZN(_01654_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05071_ (.I0(\u_cpu.rf_ram.memory[16][1] ),
    .I1(\u_cpu.rf_ram.memory[17][1] ),
    .I2(\u_cpu.rf_ram.memory[18][1] ),
    .I3(\u_cpu.rf_ram.memory[19][1] ),
    .S0(_01508_),
    .S1(_01509_),
    .Z(_01655_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05072_ (.A1(_01506_),
    .A2(_01655_),
    .B(_01519_),
    .ZN(_01656_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _05073_ (.A1(_01650_),
    .A2(_01652_),
    .B1(_01654_),
    .B2(_01656_),
    .C(_01486_),
    .ZN(_01657_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05074_ (.I0(\u_cpu.rf_ram.memory[4][1] ),
    .I1(\u_cpu.rf_ram.memory[5][1] ),
    .I2(\u_cpu.rf_ram.memory[6][1] ),
    .I3(\u_cpu.rf_ram.memory[7][1] ),
    .S0(_01523_),
    .S1(_01525_),
    .Z(_01658_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05075_ (.A1(_01493_),
    .A2(_01658_),
    .ZN(_01659_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05076_ (.I0(\u_cpu.rf_ram.memory[0][1] ),
    .I1(\u_cpu.rf_ram.memory[1][1] ),
    .I2(\u_cpu.rf_ram.memory[2][1] ),
    .I3(\u_cpu.rf_ram.memory[3][1] ),
    .S0(_01530_),
    .S1(_01532_),
    .Z(_01660_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05077_ (.A1(_01528_),
    .A2(_01660_),
    .B(_01534_),
    .ZN(_01661_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05078_ (.I0(\u_cpu.rf_ram.memory[8][1] ),
    .I1(\u_cpu.rf_ram.memory[9][1] ),
    .I2(\u_cpu.rf_ram.memory[10][1] ),
    .I3(\u_cpu.rf_ram.memory[11][1] ),
    .S0(_01523_),
    .S1(_01525_),
    .Z(_01662_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05079_ (.A1(_01528_),
    .A2(_01662_),
    .ZN(_01663_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05080_ (.I0(\u_cpu.rf_ram.memory[12][1] ),
    .I1(\u_cpu.rf_ram.memory[13][1] ),
    .I2(\u_cpu.rf_ram.memory[14][1] ),
    .I3(\u_cpu.rf_ram.memory[15][1] ),
    .S0(_01530_),
    .S1(_01532_),
    .Z(_01664_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05081_ (.A1(_01513_),
    .A2(_01664_),
    .B(_01482_),
    .ZN(_01665_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _05082_ (.A1(_01659_),
    .A2(_01661_),
    .B1(_01663_),
    .B2(_01665_),
    .C(_01541_),
    .ZN(_01666_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05083_ (.I0(\u_cpu.rf_ram.memory[36][1] ),
    .I1(\u_cpu.rf_ram.memory[37][1] ),
    .I2(\u_cpu.rf_ram.memory[38][1] ),
    .I3(\u_cpu.rf_ram.memory[39][1] ),
    .S0(_01544_),
    .S1(_01545_),
    .Z(_01667_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05084_ (.A1(_01543_),
    .A2(_01667_),
    .ZN(_01668_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05085_ (.I0(\u_cpu.rf_ram.memory[32][1] ),
    .I1(\u_cpu.rf_ram.memory[33][1] ),
    .I2(\u_cpu.rf_ram.memory[34][1] ),
    .I3(\u_cpu.rf_ram.memory[35][1] ),
    .S0(_01495_),
    .S1(_01499_),
    .Z(_01669_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05086_ (.A1(_01548_),
    .A2(_01669_),
    .B(_01518_),
    .ZN(_01670_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05087_ (.I0(\u_cpu.rf_ram.memory[40][1] ),
    .I1(\u_cpu.rf_ram.memory[41][1] ),
    .I2(\u_cpu.rf_ram.memory[42][1] ),
    .I3(\u_cpu.rf_ram.memory[43][1] ),
    .S0(_01551_),
    .S1(_01524_),
    .Z(_01671_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05088_ (.A1(_01505_),
    .A2(_01671_),
    .ZN(_01672_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05089_ (.I0(\u_cpu.rf_ram.memory[44][1] ),
    .I1(\u_cpu.rf_ram.memory[45][1] ),
    .I2(\u_cpu.rf_ram.memory[46][1] ),
    .I3(\u_cpu.rf_ram.memory[47][1] ),
    .S0(_01555_),
    .S1(_01531_),
    .Z(_01673_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05090_ (.A1(_01554_),
    .A2(_01673_),
    .B(_01558_),
    .ZN(_01674_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _05091_ (.A1(_01668_),
    .A2(_01670_),
    .B1(_01672_),
    .B2(_01674_),
    .C(_01560_),
    .ZN(_01675_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05092_ (.I0(\u_cpu.rf_ram.memory[60][1] ),
    .I1(\u_cpu.rf_ram.memory[61][1] ),
    .I2(\u_cpu.rf_ram.memory[62][1] ),
    .I3(\u_cpu.rf_ram.memory[63][1] ),
    .S0(_01562_),
    .S1(_01563_),
    .Z(_01676_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05093_ (.A1(_01464_),
    .A2(_01676_),
    .ZN(_01677_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05094_ (.I0(\u_cpu.rf_ram.memory[56][1] ),
    .I1(\u_cpu.rf_ram.memory[57][1] ),
    .I2(\u_cpu.rf_ram.memory[58][1] ),
    .I3(\u_cpu.rf_ram.memory[59][1] ),
    .S0(_01567_),
    .S1(_01568_),
    .Z(_01678_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05095_ (.A1(_01566_),
    .A2(_01678_),
    .B(_01480_),
    .ZN(_01679_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05096_ (.I0(\u_cpu.rf_ram.memory[52][1] ),
    .I1(\u_cpu.rf_ram.memory[53][1] ),
    .I2(\u_cpu.rf_ram.memory[54][1] ),
    .I3(\u_cpu.rf_ram.memory[55][1] ),
    .S0(_01572_),
    .S1(_01573_),
    .Z(_01680_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05097_ (.A1(_01571_),
    .A2(_01680_),
    .ZN(_01681_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05098_ (.I0(\u_cpu.rf_ram.memory[48][1] ),
    .I1(\u_cpu.rf_ram.memory[49][1] ),
    .I2(\u_cpu.rf_ram.memory[50][1] ),
    .I3(\u_cpu.rf_ram.memory[51][1] ),
    .S0(_01576_),
    .S1(_01577_),
    .Z(_01682_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05099_ (.A1(_01505_),
    .A2(_01682_),
    .B(_01579_),
    .ZN(_01683_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _05100_ (.A1(_01677_),
    .A2(_01679_),
    .B1(_01681_),
    .B2(_01683_),
    .C(_01581_),
    .ZN(_01684_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _05101_ (.A1(_01490_),
    .A2(_01675_),
    .A3(_01684_),
    .Z(_01685_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _05102_ (.A1(_01492_),
    .A2(_01657_),
    .A3(_01666_),
    .B(_01685_),
    .ZN(_01686_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05103_ (.I0(\u_cpu.rf_ram.memory[100][1] ),
    .I1(\u_cpu.rf_ram.memory[101][1] ),
    .I2(\u_cpu.rf_ram.memory[102][1] ),
    .I3(\u_cpu.rf_ram.memory[103][1] ),
    .S0(_01572_),
    .S1(_01573_),
    .Z(_01687_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05104_ (.A1(_01571_),
    .A2(_01687_),
    .ZN(_01688_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05105_ (.I0(\u_cpu.rf_ram.memory[96][1] ),
    .I1(\u_cpu.rf_ram.memory[97][1] ),
    .I2(\u_cpu.rf_ram.memory[98][1] ),
    .I3(\u_cpu.rf_ram.memory[99][1] ),
    .S0(_01567_),
    .S1(_01568_),
    .Z(_01689_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05106_ (.A1(_01548_),
    .A2(_01689_),
    .B(_01579_),
    .ZN(_01690_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05107_ (.I0(\u_cpu.rf_ram.memory[108][1] ),
    .I1(\u_cpu.rf_ram.memory[109][1] ),
    .I2(\u_cpu.rf_ram.memory[110][1] ),
    .I3(\u_cpu.rf_ram.memory[111][1] ),
    .S0(_01551_),
    .S1(_01524_),
    .Z(_01691_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05108_ (.A1(_01512_),
    .A2(_01691_),
    .ZN(_01692_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05109_ (.I0(\u_cpu.rf_ram.memory[104][1] ),
    .I1(\u_cpu.rf_ram.memory[105][1] ),
    .I2(\u_cpu.rf_ram.memory[106][1] ),
    .I3(\u_cpu.rf_ram.memory[107][1] ),
    .S0(_01555_),
    .S1(_01531_),
    .Z(_01693_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05110_ (.A1(_01566_),
    .A2(_01693_),
    .B(_01558_),
    .ZN(_01694_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _05111_ (.A1(_01688_),
    .A2(_01690_),
    .B1(_01692_),
    .B2(_01694_),
    .C(_01560_),
    .ZN(_01695_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05112_ (.I0(\u_cpu.rf_ram.memory[124][1] ),
    .I1(\u_cpu.rf_ram.memory[125][1] ),
    .I2(\u_cpu.rf_ram.memory[126][1] ),
    .I3(\u_cpu.rf_ram.memory[127][1] ),
    .S0(_01496_),
    .S1(_01594_),
    .Z(_01696_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05113_ (.A1(_01543_),
    .A2(_01696_),
    .ZN(_01697_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05114_ (.I0(\u_cpu.rf_ram.memory[120][1] ),
    .I1(\u_cpu.rf_ram.memory[121][1] ),
    .I2(\u_cpu.rf_ram.memory[122][1] ),
    .I3(\u_cpu.rf_ram.memory[123][1] ),
    .S0(_01598_),
    .S1(_01556_),
    .Z(_01698_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05115_ (.A1(_01597_),
    .A2(_01698_),
    .B(_01600_),
    .ZN(_01699_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05116_ (.I0(\u_cpu.rf_ram.memory[112][1] ),
    .I1(\u_cpu.rf_ram.memory[113][1] ),
    .I2(\u_cpu.rf_ram.memory[114][1] ),
    .I3(\u_cpu.rf_ram.memory[115][1] ),
    .S0(_01544_),
    .S1(_01545_),
    .Z(_01700_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05117_ (.A1(_01602_),
    .A2(_01700_),
    .ZN(_01701_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05118_ (.I0(\u_cpu.rf_ram.memory[116][1] ),
    .I1(\u_cpu.rf_ram.memory[117][1] ),
    .I2(\u_cpu.rf_ram.memory[118][1] ),
    .I3(\u_cpu.rf_ram.memory[119][1] ),
    .S0(_01576_),
    .S1(_01577_),
    .Z(_01702_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05119_ (.A1(_01554_),
    .A2(_01702_),
    .B(_01607_),
    .ZN(_01703_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _05120_ (.A1(_01697_),
    .A2(_01699_),
    .B1(_01701_),
    .B2(_01703_),
    .C(_01581_),
    .ZN(_01704_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _05121_ (.A1(_01490_),
    .A2(_01695_),
    .A3(_01704_),
    .ZN(_01705_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05122_ (.I0(\u_cpu.rf_ram.memory[92][1] ),
    .I1(\u_cpu.rf_ram.memory[93][1] ),
    .I2(\u_cpu.rf_ram.memory[94][1] ),
    .I3(\u_cpu.rf_ram.memory[95][1] ),
    .S0(_01562_),
    .S1(_01563_),
    .Z(_01706_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05123_ (.A1(_01464_),
    .A2(_01706_),
    .ZN(_01707_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05124_ (.I0(\u_cpu.rf_ram.memory[88][1] ),
    .I1(\u_cpu.rf_ram.memory[89][1] ),
    .I2(\u_cpu.rf_ram.memory[90][1] ),
    .I3(\u_cpu.rf_ram.memory[91][1] ),
    .S0(_01598_),
    .S1(_01556_),
    .Z(_01708_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05125_ (.A1(_01597_),
    .A2(_01708_),
    .B(_01600_),
    .ZN(_01709_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05126_ (.I0(\u_cpu.rf_ram.memory[80][1] ),
    .I1(\u_cpu.rf_ram.memory[81][1] ),
    .I2(\u_cpu.rf_ram.memory[82][1] ),
    .I3(\u_cpu.rf_ram.memory[83][1] ),
    .S0(_01496_),
    .S1(_01594_),
    .Z(_01710_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05127_ (.A1(_01602_),
    .A2(_01710_),
    .ZN(_01711_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05128_ (.I0(\u_cpu.rf_ram.memory[84][1] ),
    .I1(\u_cpu.rf_ram.memory[85][1] ),
    .I2(\u_cpu.rf_ram.memory[86][1] ),
    .I3(\u_cpu.rf_ram.memory[87][1] ),
    .S0(_01507_),
    .S1(_01605_),
    .Z(_01712_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05129_ (.A1(_01617_),
    .A2(_01712_),
    .B(_01607_),
    .ZN(_01713_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _05130_ (.A1(_01707_),
    .A2(_01709_),
    .B1(_01711_),
    .B2(_01713_),
    .C(_01486_),
    .ZN(_01714_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05131_ (.I0(\u_cpu.rf_ram.memory[64][1] ),
    .I1(\u_cpu.rf_ram.memory[65][1] ),
    .I2(\u_cpu.rf_ram.memory[66][1] ),
    .I3(\u_cpu.rf_ram.memory[67][1] ),
    .S0(_01522_),
    .S1(_01622_),
    .Z(_01715_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05132_ (.A1(_01621_),
    .A2(_01715_),
    .ZN(_01716_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05133_ (.I0(\u_cpu.rf_ram.memory[68][1] ),
    .I1(\u_cpu.rf_ram.memory[69][1] ),
    .I2(\u_cpu.rf_ram.memory[70][1] ),
    .I3(\u_cpu.rf_ram.memory[71][1] ),
    .S0(_01507_),
    .S1(_01605_),
    .Z(_01717_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05134_ (.A1(_01617_),
    .A2(_01717_),
    .B(_01519_),
    .ZN(_01718_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05135_ (.I0(\u_cpu.rf_ram.memory[72][1] ),
    .I1(\u_cpu.rf_ram.memory[73][1] ),
    .I2(\u_cpu.rf_ram.memory[74][1] ),
    .I3(\u_cpu.rf_ram.memory[75][1] ),
    .S0(_01522_),
    .S1(_01622_),
    .Z(_01719_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05136_ (.A1(_01621_),
    .A2(_01719_),
    .ZN(_01720_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05137_ (.I0(\u_cpu.rf_ram.memory[76][1] ),
    .I1(\u_cpu.rf_ram.memory[77][1] ),
    .I2(\u_cpu.rf_ram.memory[78][1] ),
    .I3(\u_cpu.rf_ram.memory[79][1] ),
    .S0(_01529_),
    .S1(_01500_),
    .Z(_01721_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05138_ (.A1(_01512_),
    .A2(_01721_),
    .B(_01481_),
    .ZN(_01722_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _05139_ (.A1(_01716_),
    .A2(_01718_),
    .B1(_01720_),
    .B2(_01722_),
    .C(_01541_),
    .ZN(_01723_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _05140_ (.A1(_01492_),
    .A2(_01714_),
    .A3(_01723_),
    .ZN(_01724_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05141_ (.A1(_01705_),
    .A2(_01724_),
    .B(_01471_),
    .ZN(_01725_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05142_ (.I0(\u_cpu.rf_ram.memory[128][1] ),
    .I1(\u_cpu.rf_ram.memory[129][1] ),
    .I2(\u_cpu.rf_ram.memory[130][1] ),
    .I3(\u_cpu.rf_ram.memory[131][1] ),
    .S0(_01634_),
    .S1(_01635_),
    .Z(_01726_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05143_ (.A1(_01465_),
    .A2(_01726_),
    .ZN(_01727_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05144_ (.I0(\u_cpu.rf_ram.memory[132][1] ),
    .I1(\u_cpu.rf_ram.memory[133][1] ),
    .I2(\u_cpu.rf_ram.memory[134][1] ),
    .I3(\u_cpu.rf_ram.memory[135][1] ),
    .S0(_01634_),
    .S1(_01635_),
    .Z(_01728_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05145_ (.A1(_01638_),
    .A2(_01728_),
    .B(_01482_),
    .ZN(_01729_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05146_ (.I0(\u_cpu.rf_ram.memory[136][1] ),
    .I1(\u_cpu.rf_ram.memory[137][1] ),
    .I2(\u_cpu.rf_ram.memory[138][1] ),
    .I3(\u_cpu.rf_ram.memory[139][1] ),
    .S0(_01641_),
    .S1(_01642_),
    .Z(_01730_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05147_ (.A1(_01465_),
    .A2(_01730_),
    .ZN(_01731_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05148_ (.I0(\u_cpu.rf_ram.memory[140][1] ),
    .I1(\u_cpu.rf_ram.memory[141][1] ),
    .I2(\u_cpu.rf_ram.memory[142][1] ),
    .I3(\u_cpu.rf_ram.memory[143][1] ),
    .S0(_01641_),
    .S1(_01642_),
    .Z(_01732_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05149_ (.A1(_01638_),
    .A2(_01732_),
    .B(_01534_),
    .ZN(_01733_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _05150_ (.A1(_01727_),
    .A2(_01729_),
    .B1(_01731_),
    .B2(_01733_),
    .C(_01466_),
    .ZN(_01734_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05151_ (.A1(_01725_),
    .A2(_01734_),
    .ZN(_01735_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05152_ (.A1(_01473_),
    .A2(_01686_),
    .B(_01735_),
    .ZN(_00001_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05153_ (.I0(\u_cpu.rf_ram.memory[28][2] ),
    .I1(\u_cpu.rf_ram.memory[29][2] ),
    .I2(\u_cpu.rf_ram.memory[30][2] ),
    .I3(\u_cpu.rf_ram.memory[31][2] ),
    .S0(_01497_),
    .S1(_01501_),
    .Z(_01736_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05154_ (.A1(_01493_),
    .A2(_01736_),
    .ZN(_01737_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05155_ (.I0(\u_cpu.rf_ram.memory[24][2] ),
    .I1(\u_cpu.rf_ram.memory[25][2] ),
    .I2(\u_cpu.rf_ram.memory[26][2] ),
    .I3(\u_cpu.rf_ram.memory[27][2] ),
    .S0(_01508_),
    .S1(_01509_),
    .Z(_01738_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05156_ (.A1(_01506_),
    .A2(_01738_),
    .B(_01481_),
    .ZN(_01739_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05157_ (.I0(\u_cpu.rf_ram.memory[20][2] ),
    .I1(\u_cpu.rf_ram.memory[21][2] ),
    .I2(\u_cpu.rf_ram.memory[22][2] ),
    .I3(\u_cpu.rf_ram.memory[23][2] ),
    .S0(_01497_),
    .S1(_01501_),
    .Z(_01740_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05158_ (.A1(_01513_),
    .A2(_01740_),
    .ZN(_01741_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05159_ (.I0(\u_cpu.rf_ram.memory[16][2] ),
    .I1(\u_cpu.rf_ram.memory[17][2] ),
    .I2(\u_cpu.rf_ram.memory[18][2] ),
    .I3(\u_cpu.rf_ram.memory[19][2] ),
    .S0(_01508_),
    .S1(_01509_),
    .Z(_01742_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05160_ (.A1(_01506_),
    .A2(_01742_),
    .B(_01519_),
    .ZN(_01743_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _05161_ (.A1(_01737_),
    .A2(_01739_),
    .B1(_01741_),
    .B2(_01743_),
    .C(_01486_),
    .ZN(_01744_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05162_ (.I0(\u_cpu.rf_ram.memory[4][2] ),
    .I1(\u_cpu.rf_ram.memory[5][2] ),
    .I2(\u_cpu.rf_ram.memory[6][2] ),
    .I3(\u_cpu.rf_ram.memory[7][2] ),
    .S0(_01523_),
    .S1(_01525_),
    .Z(_01745_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05163_ (.A1(_01493_),
    .A2(_01745_),
    .ZN(_01746_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05164_ (.I0(\u_cpu.rf_ram.memory[0][2] ),
    .I1(\u_cpu.rf_ram.memory[1][2] ),
    .I2(\u_cpu.rf_ram.memory[2][2] ),
    .I3(\u_cpu.rf_ram.memory[3][2] ),
    .S0(_01530_),
    .S1(_01532_),
    .Z(_01747_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05165_ (.A1(_01528_),
    .A2(_01747_),
    .B(_01534_),
    .ZN(_01748_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05166_ (.I0(\u_cpu.rf_ram.memory[8][2] ),
    .I1(\u_cpu.rf_ram.memory[9][2] ),
    .I2(\u_cpu.rf_ram.memory[10][2] ),
    .I3(\u_cpu.rf_ram.memory[11][2] ),
    .S0(_01523_),
    .S1(_01525_),
    .Z(_01749_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05167_ (.A1(_01528_),
    .A2(_01749_),
    .ZN(_01750_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05168_ (.I0(\u_cpu.rf_ram.memory[12][2] ),
    .I1(\u_cpu.rf_ram.memory[13][2] ),
    .I2(\u_cpu.rf_ram.memory[14][2] ),
    .I3(\u_cpu.rf_ram.memory[15][2] ),
    .S0(_01530_),
    .S1(_01532_),
    .Z(_01751_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05169_ (.A1(_01513_),
    .A2(_01751_),
    .B(_01482_),
    .ZN(_01752_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _05170_ (.A1(_01746_),
    .A2(_01748_),
    .B1(_01750_),
    .B2(_01752_),
    .C(_01541_),
    .ZN(_01753_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05171_ (.I0(\u_cpu.rf_ram.memory[36][2] ),
    .I1(\u_cpu.rf_ram.memory[37][2] ),
    .I2(\u_cpu.rf_ram.memory[38][2] ),
    .I3(\u_cpu.rf_ram.memory[39][2] ),
    .S0(_01544_),
    .S1(_01545_),
    .Z(_01754_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05172_ (.A1(_01543_),
    .A2(_01754_),
    .ZN(_01755_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05173_ (.I0(\u_cpu.rf_ram.memory[32][2] ),
    .I1(\u_cpu.rf_ram.memory[33][2] ),
    .I2(\u_cpu.rf_ram.memory[34][2] ),
    .I3(\u_cpu.rf_ram.memory[35][2] ),
    .S0(_01495_),
    .S1(_01499_),
    .Z(_01756_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05174_ (.A1(_01548_),
    .A2(_01756_),
    .B(_01518_),
    .ZN(_01757_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05175_ (.I0(\u_cpu.rf_ram.memory[40][2] ),
    .I1(\u_cpu.rf_ram.memory[41][2] ),
    .I2(\u_cpu.rf_ram.memory[42][2] ),
    .I3(\u_cpu.rf_ram.memory[43][2] ),
    .S0(_01551_),
    .S1(_01524_),
    .Z(_01758_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05176_ (.A1(_01505_),
    .A2(_01758_),
    .ZN(_01759_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05177_ (.I0(\u_cpu.rf_ram.memory[44][2] ),
    .I1(\u_cpu.rf_ram.memory[45][2] ),
    .I2(\u_cpu.rf_ram.memory[46][2] ),
    .I3(\u_cpu.rf_ram.memory[47][2] ),
    .S0(_01555_),
    .S1(_01531_),
    .Z(_01760_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05178_ (.A1(_01554_),
    .A2(_01760_),
    .B(_01558_),
    .ZN(_01761_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _05179_ (.A1(_01755_),
    .A2(_01757_),
    .B1(_01759_),
    .B2(_01761_),
    .C(_01560_),
    .ZN(_01762_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05180_ (.I0(\u_cpu.rf_ram.memory[60][2] ),
    .I1(\u_cpu.rf_ram.memory[61][2] ),
    .I2(\u_cpu.rf_ram.memory[62][2] ),
    .I3(\u_cpu.rf_ram.memory[63][2] ),
    .S0(_01562_),
    .S1(_01563_),
    .Z(_01763_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05181_ (.A1(_01464_),
    .A2(_01763_),
    .ZN(_01764_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05182_ (.I0(\u_cpu.rf_ram.memory[56][2] ),
    .I1(\u_cpu.rf_ram.memory[57][2] ),
    .I2(\u_cpu.rf_ram.memory[58][2] ),
    .I3(\u_cpu.rf_ram.memory[59][2] ),
    .S0(_01567_),
    .S1(_01568_),
    .Z(_01765_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05183_ (.A1(_01566_),
    .A2(_01765_),
    .B(_01480_),
    .ZN(_01766_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05184_ (.I0(\u_cpu.rf_ram.memory[52][2] ),
    .I1(\u_cpu.rf_ram.memory[53][2] ),
    .I2(\u_cpu.rf_ram.memory[54][2] ),
    .I3(\u_cpu.rf_ram.memory[55][2] ),
    .S0(_01572_),
    .S1(_01573_),
    .Z(_01767_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05185_ (.A1(_01571_),
    .A2(_01767_),
    .ZN(_01768_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05186_ (.I0(\u_cpu.rf_ram.memory[48][2] ),
    .I1(\u_cpu.rf_ram.memory[49][2] ),
    .I2(\u_cpu.rf_ram.memory[50][2] ),
    .I3(\u_cpu.rf_ram.memory[51][2] ),
    .S0(_01576_),
    .S1(_01577_),
    .Z(_01769_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05187_ (.A1(_01505_),
    .A2(_01769_),
    .B(_01579_),
    .ZN(_01770_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _05188_ (.A1(_01764_),
    .A2(_01766_),
    .B1(_01768_),
    .B2(_01770_),
    .C(_01581_),
    .ZN(_01771_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _05189_ (.A1(_01490_),
    .A2(_01762_),
    .A3(_01771_),
    .Z(_01772_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _05190_ (.A1(_01492_),
    .A2(_01744_),
    .A3(_01753_),
    .B(_01772_),
    .ZN(_01773_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05191_ (.I0(\u_cpu.rf_ram.memory[100][2] ),
    .I1(\u_cpu.rf_ram.memory[101][2] ),
    .I2(\u_cpu.rf_ram.memory[102][2] ),
    .I3(\u_cpu.rf_ram.memory[103][2] ),
    .S0(_01551_),
    .S1(_01573_),
    .Z(_01774_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05192_ (.A1(_01571_),
    .A2(_01774_),
    .ZN(_01775_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05193_ (.I0(\u_cpu.rf_ram.memory[96][2] ),
    .I1(\u_cpu.rf_ram.memory[97][2] ),
    .I2(\u_cpu.rf_ram.memory[98][2] ),
    .I3(\u_cpu.rf_ram.memory[99][2] ),
    .S0(_01567_),
    .S1(_01568_),
    .Z(_01776_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05194_ (.A1(_01548_),
    .A2(_01776_),
    .B(_01579_),
    .ZN(_01777_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05195_ (.I0(\u_cpu.rf_ram.memory[108][2] ),
    .I1(\u_cpu.rf_ram.memory[109][2] ),
    .I2(\u_cpu.rf_ram.memory[110][2] ),
    .I3(\u_cpu.rf_ram.memory[111][2] ),
    .S0(_01529_),
    .S1(_01524_),
    .Z(_01778_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05196_ (.A1(_01512_),
    .A2(_01778_),
    .ZN(_01779_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05197_ (.I0(\u_cpu.rf_ram.memory[104][2] ),
    .I1(\u_cpu.rf_ram.memory[105][2] ),
    .I2(\u_cpu.rf_ram.memory[106][2] ),
    .I3(\u_cpu.rf_ram.memory[107][2] ),
    .S0(_01555_),
    .S1(_01531_),
    .Z(_01780_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05198_ (.A1(_01566_),
    .A2(_01780_),
    .B(_01558_),
    .ZN(_01781_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _05199_ (.A1(_01775_),
    .A2(_01777_),
    .B1(_01779_),
    .B2(_01781_),
    .C(_01560_),
    .ZN(_01782_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05200_ (.I0(\u_cpu.rf_ram.memory[124][2] ),
    .I1(\u_cpu.rf_ram.memory[125][2] ),
    .I2(\u_cpu.rf_ram.memory[126][2] ),
    .I3(\u_cpu.rf_ram.memory[127][2] ),
    .S0(_01496_),
    .S1(_01594_),
    .Z(_01783_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05201_ (.A1(_01543_),
    .A2(_01783_),
    .ZN(_01784_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05202_ (.I0(\u_cpu.rf_ram.memory[120][2] ),
    .I1(\u_cpu.rf_ram.memory[121][2] ),
    .I2(\u_cpu.rf_ram.memory[122][2] ),
    .I3(\u_cpu.rf_ram.memory[123][2] ),
    .S0(_01598_),
    .S1(_01556_),
    .Z(_01785_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05203_ (.A1(_01597_),
    .A2(_01785_),
    .B(_01600_),
    .ZN(_01786_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05204_ (.I0(\u_cpu.rf_ram.memory[112][2] ),
    .I1(\u_cpu.rf_ram.memory[113][2] ),
    .I2(\u_cpu.rf_ram.memory[114][2] ),
    .I3(\u_cpu.rf_ram.memory[115][2] ),
    .S0(_01572_),
    .S1(_01545_),
    .Z(_01787_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05205_ (.A1(_01602_),
    .A2(_01787_),
    .ZN(_01788_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05206_ (.I0(\u_cpu.rf_ram.memory[116][2] ),
    .I1(\u_cpu.rf_ram.memory[117][2] ),
    .I2(\u_cpu.rf_ram.memory[118][2] ),
    .I3(\u_cpu.rf_ram.memory[119][2] ),
    .S0(_01576_),
    .S1(_01577_),
    .Z(_01789_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05207_ (.A1(_01554_),
    .A2(_01789_),
    .B(_01607_),
    .ZN(_01790_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _05208_ (.A1(_01784_),
    .A2(_01786_),
    .B1(_01788_),
    .B2(_01790_),
    .C(_01581_),
    .ZN(_01791_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _05209_ (.A1(_01490_),
    .A2(_01782_),
    .A3(_01791_),
    .ZN(_01792_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05210_ (.I0(\u_cpu.rf_ram.memory[92][2] ),
    .I1(\u_cpu.rf_ram.memory[93][2] ),
    .I2(\u_cpu.rf_ram.memory[94][2] ),
    .I3(\u_cpu.rf_ram.memory[95][2] ),
    .S0(_01562_),
    .S1(_01563_),
    .Z(_01793_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05211_ (.A1(_01464_),
    .A2(_01793_),
    .ZN(_01794_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05212_ (.I0(\u_cpu.rf_ram.memory[88][2] ),
    .I1(\u_cpu.rf_ram.memory[89][2] ),
    .I2(\u_cpu.rf_ram.memory[90][2] ),
    .I3(\u_cpu.rf_ram.memory[91][2] ),
    .S0(_01598_),
    .S1(_01556_),
    .Z(_01795_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05213_ (.A1(_01597_),
    .A2(_01795_),
    .B(_01600_),
    .ZN(_01796_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05214_ (.I0(\u_cpu.rf_ram.memory[80][2] ),
    .I1(\u_cpu.rf_ram.memory[81][2] ),
    .I2(\u_cpu.rf_ram.memory[82][2] ),
    .I3(\u_cpu.rf_ram.memory[83][2] ),
    .S0(_01544_),
    .S1(_01594_),
    .Z(_01797_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05215_ (.A1(_01602_),
    .A2(_01797_),
    .ZN(_01798_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05216_ (.I0(\u_cpu.rf_ram.memory[84][2] ),
    .I1(\u_cpu.rf_ram.memory[85][2] ),
    .I2(\u_cpu.rf_ram.memory[86][2] ),
    .I3(\u_cpu.rf_ram.memory[87][2] ),
    .S0(_01507_),
    .S1(_01605_),
    .Z(_01799_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05217_ (.A1(_01617_),
    .A2(_01799_),
    .B(_01607_),
    .ZN(_01800_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _05218_ (.A1(_01794_),
    .A2(_01796_),
    .B1(_01798_),
    .B2(_01800_),
    .C(_01486_),
    .ZN(_01801_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05219_ (.I0(\u_cpu.rf_ram.memory[64][2] ),
    .I1(\u_cpu.rf_ram.memory[65][2] ),
    .I2(\u_cpu.rf_ram.memory[66][2] ),
    .I3(\u_cpu.rf_ram.memory[67][2] ),
    .S0(_01522_),
    .S1(_01622_),
    .Z(_01802_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05220_ (.A1(_01621_),
    .A2(_01802_),
    .ZN(_01803_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05221_ (.I0(\u_cpu.rf_ram.memory[68][2] ),
    .I1(\u_cpu.rf_ram.memory[69][2] ),
    .I2(\u_cpu.rf_ram.memory[70][2] ),
    .I3(\u_cpu.rf_ram.memory[71][2] ),
    .S0(_01507_),
    .S1(_01605_),
    .Z(_01804_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05222_ (.A1(_01617_),
    .A2(_01804_),
    .B(_01519_),
    .ZN(_01805_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05223_ (.I0(\u_cpu.rf_ram.memory[72][2] ),
    .I1(\u_cpu.rf_ram.memory[73][2] ),
    .I2(\u_cpu.rf_ram.memory[74][2] ),
    .I3(\u_cpu.rf_ram.memory[75][2] ),
    .S0(_01522_),
    .S1(_01622_),
    .Z(_01806_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05224_ (.A1(_01621_),
    .A2(_01806_),
    .ZN(_01807_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05225_ (.I0(\u_cpu.rf_ram.memory[76][2] ),
    .I1(\u_cpu.rf_ram.memory[77][2] ),
    .I2(\u_cpu.rf_ram.memory[78][2] ),
    .I3(\u_cpu.rf_ram.memory[79][2] ),
    .S0(_01529_),
    .S1(_01500_),
    .Z(_01808_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05226_ (.A1(_01512_),
    .A2(_01808_),
    .B(_01481_),
    .ZN(_01809_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _05227_ (.A1(_01803_),
    .A2(_01805_),
    .B1(_01807_),
    .B2(_01809_),
    .C(_01541_),
    .ZN(_01810_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _05228_ (.A1(_01492_),
    .A2(_01801_),
    .A3(_01810_),
    .ZN(_01811_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05229_ (.A1(_01792_),
    .A2(_01811_),
    .B(_01471_),
    .ZN(_01812_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05230_ (.I0(\u_cpu.rf_ram.memory[136][2] ),
    .I1(\u_cpu.rf_ram.memory[137][2] ),
    .I2(\u_cpu.rf_ram.memory[138][2] ),
    .I3(\u_cpu.rf_ram.memory[139][2] ),
    .S0(_01634_),
    .S1(_01635_),
    .Z(_01813_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05231_ (.A1(_01465_),
    .A2(_01813_),
    .ZN(_01814_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05232_ (.I0(\u_cpu.rf_ram.memory[140][2] ),
    .I1(\u_cpu.rf_ram.memory[141][2] ),
    .I2(\u_cpu.rf_ram.memory[142][2] ),
    .I3(\u_cpu.rf_ram.memory[143][2] ),
    .S0(_01634_),
    .S1(_01635_),
    .Z(_01815_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05233_ (.A1(_01638_),
    .A2(_01815_),
    .B(_01534_),
    .ZN(_01816_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05234_ (.I0(\u_cpu.rf_ram.memory[128][2] ),
    .I1(\u_cpu.rf_ram.memory[129][2] ),
    .I2(\u_cpu.rf_ram.memory[130][2] ),
    .I3(\u_cpu.rf_ram.memory[131][2] ),
    .S0(_01641_),
    .S1(_01642_),
    .Z(_01817_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05235_ (.A1(_01465_),
    .A2(_01817_),
    .ZN(_01818_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05236_ (.I0(\u_cpu.rf_ram.memory[132][2] ),
    .I1(\u_cpu.rf_ram.memory[133][2] ),
    .I2(\u_cpu.rf_ram.memory[134][2] ),
    .I3(\u_cpu.rf_ram.memory[135][2] ),
    .S0(_01641_),
    .S1(_01642_),
    .Z(_01819_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05237_ (.A1(_01638_),
    .A2(_01819_),
    .B(_01482_),
    .ZN(_01820_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _05238_ (.A1(_01814_),
    .A2(_01816_),
    .B1(_01818_),
    .B2(_01820_),
    .C(_01466_),
    .ZN(_01821_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05239_ (.A1(_01812_),
    .A2(_01821_),
    .ZN(_01822_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05240_ (.A1(_01473_),
    .A2(_01773_),
    .B(_01822_),
    .ZN(_00002_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05241_ (.I0(\u_cpu.rf_ram.memory[28][3] ),
    .I1(\u_cpu.rf_ram.memory[29][3] ),
    .I2(\u_cpu.rf_ram.memory[30][3] ),
    .I3(\u_cpu.rf_ram.memory[31][3] ),
    .S0(_01497_),
    .S1(_01501_),
    .Z(_01823_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05242_ (.A1(_01493_),
    .A2(_01823_),
    .ZN(_01824_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05243_ (.I0(\u_cpu.rf_ram.memory[24][3] ),
    .I1(\u_cpu.rf_ram.memory[25][3] ),
    .I2(\u_cpu.rf_ram.memory[26][3] ),
    .I3(\u_cpu.rf_ram.memory[27][3] ),
    .S0(_01508_),
    .S1(_01509_),
    .Z(_01825_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05244_ (.A1(_01506_),
    .A2(_01825_),
    .B(_01481_),
    .ZN(_01826_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05245_ (.I0(\u_cpu.rf_ram.memory[20][3] ),
    .I1(\u_cpu.rf_ram.memory[21][3] ),
    .I2(\u_cpu.rf_ram.memory[22][3] ),
    .I3(\u_cpu.rf_ram.memory[23][3] ),
    .S0(_01497_),
    .S1(_01501_),
    .Z(_01827_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05246_ (.A1(_01513_),
    .A2(_01827_),
    .ZN(_01828_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05247_ (.I0(\u_cpu.rf_ram.memory[16][3] ),
    .I1(\u_cpu.rf_ram.memory[17][3] ),
    .I2(\u_cpu.rf_ram.memory[18][3] ),
    .I3(\u_cpu.rf_ram.memory[19][3] ),
    .S0(_01508_),
    .S1(_01509_),
    .Z(_01829_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05248_ (.A1(_01506_),
    .A2(_01829_),
    .B(_01519_),
    .ZN(_01830_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _05249_ (.A1(_01824_),
    .A2(_01826_),
    .B1(_01828_),
    .B2(_01830_),
    .C(_01486_),
    .ZN(_01831_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05250_ (.I0(\u_cpu.rf_ram.memory[4][3] ),
    .I1(\u_cpu.rf_ram.memory[5][3] ),
    .I2(\u_cpu.rf_ram.memory[6][3] ),
    .I3(\u_cpu.rf_ram.memory[7][3] ),
    .S0(_01523_),
    .S1(_01525_),
    .Z(_01832_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05251_ (.A1(_01493_),
    .A2(_01832_),
    .ZN(_01833_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05252_ (.I0(\u_cpu.rf_ram.memory[0][3] ),
    .I1(\u_cpu.rf_ram.memory[1][3] ),
    .I2(\u_cpu.rf_ram.memory[2][3] ),
    .I3(\u_cpu.rf_ram.memory[3][3] ),
    .S0(_01530_),
    .S1(_01532_),
    .Z(_01834_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05253_ (.A1(_01528_),
    .A2(_01834_),
    .B(_01534_),
    .ZN(_01835_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05254_ (.I0(\u_cpu.rf_ram.memory[8][3] ),
    .I1(\u_cpu.rf_ram.memory[9][3] ),
    .I2(\u_cpu.rf_ram.memory[10][3] ),
    .I3(\u_cpu.rf_ram.memory[11][3] ),
    .S0(_01523_),
    .S1(_01525_),
    .Z(_01836_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05255_ (.A1(_01528_),
    .A2(_01836_),
    .ZN(_01837_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05256_ (.I0(\u_cpu.rf_ram.memory[12][3] ),
    .I1(\u_cpu.rf_ram.memory[13][3] ),
    .I2(\u_cpu.rf_ram.memory[14][3] ),
    .I3(\u_cpu.rf_ram.memory[15][3] ),
    .S0(_01530_),
    .S1(_01532_),
    .Z(_01838_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05257_ (.A1(_01513_),
    .A2(_01838_),
    .B(_01482_),
    .ZN(_01839_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _05258_ (.A1(_01833_),
    .A2(_01835_),
    .B1(_01837_),
    .B2(_01839_),
    .C(_01541_),
    .ZN(_01840_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05259_ (.I0(\u_cpu.rf_ram.memory[36][3] ),
    .I1(\u_cpu.rf_ram.memory[37][3] ),
    .I2(\u_cpu.rf_ram.memory[38][3] ),
    .I3(\u_cpu.rf_ram.memory[39][3] ),
    .S0(_01544_),
    .S1(_01545_),
    .Z(_01841_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05260_ (.A1(_01543_),
    .A2(_01841_),
    .ZN(_01842_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05261_ (.I0(\u_cpu.rf_ram.memory[32][3] ),
    .I1(\u_cpu.rf_ram.memory[33][3] ),
    .I2(\u_cpu.rf_ram.memory[34][3] ),
    .I3(\u_cpu.rf_ram.memory[35][3] ),
    .S0(_01495_),
    .S1(_01499_),
    .Z(_01843_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05262_ (.A1(_01548_),
    .A2(_01843_),
    .B(_01518_),
    .ZN(_01844_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05263_ (.I0(\u_cpu.rf_ram.memory[40][3] ),
    .I1(\u_cpu.rf_ram.memory[41][3] ),
    .I2(\u_cpu.rf_ram.memory[42][3] ),
    .I3(\u_cpu.rf_ram.memory[43][3] ),
    .S0(_01551_),
    .S1(_01524_),
    .Z(_01845_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05264_ (.A1(_01505_),
    .A2(_01845_),
    .ZN(_01846_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05265_ (.I0(\u_cpu.rf_ram.memory[44][3] ),
    .I1(\u_cpu.rf_ram.memory[45][3] ),
    .I2(\u_cpu.rf_ram.memory[46][3] ),
    .I3(\u_cpu.rf_ram.memory[47][3] ),
    .S0(_01555_),
    .S1(_01531_),
    .Z(_01847_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05266_ (.A1(_01554_),
    .A2(_01847_),
    .B(_01558_),
    .ZN(_01848_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _05267_ (.A1(_01842_),
    .A2(_01844_),
    .B1(_01846_),
    .B2(_01848_),
    .C(_01560_),
    .ZN(_01849_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05268_ (.I0(\u_cpu.rf_ram.memory[60][3] ),
    .I1(\u_cpu.rf_ram.memory[61][3] ),
    .I2(\u_cpu.rf_ram.memory[62][3] ),
    .I3(\u_cpu.rf_ram.memory[63][3] ),
    .S0(_01496_),
    .S1(_01563_),
    .Z(_01850_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05269_ (.A1(_01464_),
    .A2(_01850_),
    .ZN(_01851_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05270_ (.I0(\u_cpu.rf_ram.memory[56][3] ),
    .I1(\u_cpu.rf_ram.memory[57][3] ),
    .I2(\u_cpu.rf_ram.memory[58][3] ),
    .I3(\u_cpu.rf_ram.memory[59][3] ),
    .S0(_01567_),
    .S1(_01568_),
    .Z(_01852_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05271_ (.A1(_01566_),
    .A2(_01852_),
    .B(_01480_),
    .ZN(_01853_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05272_ (.I0(\u_cpu.rf_ram.memory[52][3] ),
    .I1(\u_cpu.rf_ram.memory[53][3] ),
    .I2(\u_cpu.rf_ram.memory[54][3] ),
    .I3(\u_cpu.rf_ram.memory[55][3] ),
    .S0(_01572_),
    .S1(_01573_),
    .Z(_01854_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05273_ (.A1(_01571_),
    .A2(_01854_),
    .ZN(_01855_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05274_ (.I0(\u_cpu.rf_ram.memory[48][3] ),
    .I1(\u_cpu.rf_ram.memory[49][3] ),
    .I2(\u_cpu.rf_ram.memory[50][3] ),
    .I3(\u_cpu.rf_ram.memory[51][3] ),
    .S0(_01576_),
    .S1(_01577_),
    .Z(_01856_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05275_ (.A1(_01505_),
    .A2(_01856_),
    .B(_01579_),
    .ZN(_01857_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _05276_ (.A1(_01851_),
    .A2(_01853_),
    .B1(_01855_),
    .B2(_01857_),
    .C(_01581_),
    .ZN(_01858_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _05277_ (.A1(_01490_),
    .A2(_01849_),
    .A3(_01858_),
    .Z(_01859_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _05278_ (.A1(_01492_),
    .A2(_01831_),
    .A3(_01840_),
    .B(_01859_),
    .ZN(_01860_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05279_ (.I0(\u_cpu.rf_ram.memory[100][3] ),
    .I1(\u_cpu.rf_ram.memory[101][3] ),
    .I2(\u_cpu.rf_ram.memory[102][3] ),
    .I3(\u_cpu.rf_ram.memory[103][3] ),
    .S0(_01551_),
    .S1(_01573_),
    .Z(_01861_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05280_ (.A1(_01571_),
    .A2(_01861_),
    .ZN(_01862_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05281_ (.I0(\u_cpu.rf_ram.memory[96][3] ),
    .I1(\u_cpu.rf_ram.memory[97][3] ),
    .I2(\u_cpu.rf_ram.memory[98][3] ),
    .I3(\u_cpu.rf_ram.memory[99][3] ),
    .S0(_01567_),
    .S1(_01568_),
    .Z(_01863_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05282_ (.A1(_01548_),
    .A2(_01863_),
    .B(_01579_),
    .ZN(_01864_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05283_ (.I0(\u_cpu.rf_ram.memory[108][3] ),
    .I1(\u_cpu.rf_ram.memory[109][3] ),
    .I2(\u_cpu.rf_ram.memory[110][3] ),
    .I3(\u_cpu.rf_ram.memory[111][3] ),
    .S0(_01529_),
    .S1(_01500_),
    .Z(_01865_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05284_ (.A1(_01512_),
    .A2(_01865_),
    .ZN(_01866_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05285_ (.I0(\u_cpu.rf_ram.memory[104][3] ),
    .I1(\u_cpu.rf_ram.memory[105][3] ),
    .I2(\u_cpu.rf_ram.memory[106][3] ),
    .I3(\u_cpu.rf_ram.memory[107][3] ),
    .S0(_01555_),
    .S1(_01531_),
    .Z(_01867_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05286_ (.A1(_01566_),
    .A2(_01867_),
    .B(_01558_),
    .ZN(_01868_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _05287_ (.A1(_01862_),
    .A2(_01864_),
    .B1(_01866_),
    .B2(_01868_),
    .C(_01560_),
    .ZN(_01869_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05288_ (.I0(\u_cpu.rf_ram.memory[124][3] ),
    .I1(\u_cpu.rf_ram.memory[125][3] ),
    .I2(\u_cpu.rf_ram.memory[126][3] ),
    .I3(\u_cpu.rf_ram.memory[127][3] ),
    .S0(_01496_),
    .S1(_01594_),
    .Z(_01870_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05289_ (.A1(_01543_),
    .A2(_01870_),
    .ZN(_01871_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05290_ (.I0(\u_cpu.rf_ram.memory[120][3] ),
    .I1(\u_cpu.rf_ram.memory[121][3] ),
    .I2(\u_cpu.rf_ram.memory[122][3] ),
    .I3(\u_cpu.rf_ram.memory[123][3] ),
    .S0(_01598_),
    .S1(_01556_),
    .Z(_01872_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05291_ (.A1(_01597_),
    .A2(_01872_),
    .B(_01600_),
    .ZN(_01873_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05292_ (.I0(\u_cpu.rf_ram.memory[112][3] ),
    .I1(\u_cpu.rf_ram.memory[113][3] ),
    .I2(\u_cpu.rf_ram.memory[114][3] ),
    .I3(\u_cpu.rf_ram.memory[115][3] ),
    .S0(_01572_),
    .S1(_01545_),
    .Z(_01874_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05293_ (.A1(_01602_),
    .A2(_01874_),
    .ZN(_01875_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05294_ (.I0(\u_cpu.rf_ram.memory[116][3] ),
    .I1(\u_cpu.rf_ram.memory[117][3] ),
    .I2(\u_cpu.rf_ram.memory[118][3] ),
    .I3(\u_cpu.rf_ram.memory[119][3] ),
    .S0(_01576_),
    .S1(_01577_),
    .Z(_01876_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05295_ (.A1(_01554_),
    .A2(_01876_),
    .B(_01607_),
    .ZN(_01877_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _05296_ (.A1(_01871_),
    .A2(_01873_),
    .B1(_01875_),
    .B2(_01877_),
    .C(_01581_),
    .ZN(_01878_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _05297_ (.A1(_01490_),
    .A2(_01869_),
    .A3(_01878_),
    .ZN(_01879_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05298_ (.I0(\u_cpu.rf_ram.memory[92][3] ),
    .I1(\u_cpu.rf_ram.memory[93][3] ),
    .I2(\u_cpu.rf_ram.memory[94][3] ),
    .I3(\u_cpu.rf_ram.memory[95][3] ),
    .S0(_01562_),
    .S1(_01563_),
    .Z(_01880_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05299_ (.A1(_01464_),
    .A2(_01880_),
    .ZN(_01881_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05300_ (.I0(\u_cpu.rf_ram.memory[88][3] ),
    .I1(\u_cpu.rf_ram.memory[89][3] ),
    .I2(\u_cpu.rf_ram.memory[90][3] ),
    .I3(\u_cpu.rf_ram.memory[91][3] ),
    .S0(_01598_),
    .S1(_01556_),
    .Z(_01882_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05301_ (.A1(_01597_),
    .A2(_01882_),
    .B(_01600_),
    .ZN(_01883_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05302_ (.I0(\u_cpu.rf_ram.memory[80][3] ),
    .I1(\u_cpu.rf_ram.memory[81][3] ),
    .I2(\u_cpu.rf_ram.memory[82][3] ),
    .I3(\u_cpu.rf_ram.memory[83][3] ),
    .S0(_01544_),
    .S1(_01594_),
    .Z(_01884_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05303_ (.A1(_01602_),
    .A2(_01884_),
    .ZN(_01885_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05304_ (.I0(\u_cpu.rf_ram.memory[84][3] ),
    .I1(\u_cpu.rf_ram.memory[85][3] ),
    .I2(\u_cpu.rf_ram.memory[86][3] ),
    .I3(\u_cpu.rf_ram.memory[87][3] ),
    .S0(_01507_),
    .S1(_01605_),
    .Z(_01886_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05305_ (.A1(_01617_),
    .A2(_01886_),
    .B(_01607_),
    .ZN(_01887_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _05306_ (.A1(_01881_),
    .A2(_01883_),
    .B1(_01885_),
    .B2(_01887_),
    .C(_01486_),
    .ZN(_01888_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05307_ (.I0(\u_cpu.rf_ram.memory[64][3] ),
    .I1(\u_cpu.rf_ram.memory[65][3] ),
    .I2(\u_cpu.rf_ram.memory[66][3] ),
    .I3(\u_cpu.rf_ram.memory[67][3] ),
    .S0(_01522_),
    .S1(_01622_),
    .Z(_01889_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05308_ (.A1(_01621_),
    .A2(_01889_),
    .ZN(_01890_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05309_ (.I0(\u_cpu.rf_ram.memory[68][3] ),
    .I1(\u_cpu.rf_ram.memory[69][3] ),
    .I2(\u_cpu.rf_ram.memory[70][3] ),
    .I3(\u_cpu.rf_ram.memory[71][3] ),
    .S0(_01507_),
    .S1(_01605_),
    .Z(_01891_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05310_ (.A1(_01617_),
    .A2(_01891_),
    .B(_01519_),
    .ZN(_01892_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05311_ (.I0(\u_cpu.rf_ram.memory[72][3] ),
    .I1(\u_cpu.rf_ram.memory[73][3] ),
    .I2(\u_cpu.rf_ram.memory[74][3] ),
    .I3(\u_cpu.rf_ram.memory[75][3] ),
    .S0(_01562_),
    .S1(_01622_),
    .Z(_01893_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05312_ (.A1(_01621_),
    .A2(_01893_),
    .ZN(_01894_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05313_ (.I0(\u_cpu.rf_ram.memory[76][3] ),
    .I1(\u_cpu.rf_ram.memory[77][3] ),
    .I2(\u_cpu.rf_ram.memory[78][3] ),
    .I3(\u_cpu.rf_ram.memory[79][3] ),
    .S0(_01529_),
    .S1(_01500_),
    .Z(_01895_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05314_ (.A1(_01512_),
    .A2(_01895_),
    .B(_01481_),
    .ZN(_01896_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _05315_ (.A1(_01890_),
    .A2(_01892_),
    .B1(_01894_),
    .B2(_01896_),
    .C(_01541_),
    .ZN(_01897_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _05316_ (.A1(_01492_),
    .A2(_01888_),
    .A3(_01897_),
    .ZN(_01898_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05317_ (.A1(_01879_),
    .A2(_01898_),
    .B(_01471_),
    .ZN(_01899_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05318_ (.I0(\u_cpu.rf_ram.memory[128][3] ),
    .I1(\u_cpu.rf_ram.memory[129][3] ),
    .I2(\u_cpu.rf_ram.memory[130][3] ),
    .I3(\u_cpu.rf_ram.memory[131][3] ),
    .S0(_01634_),
    .S1(_01635_),
    .Z(_01900_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05319_ (.A1(_01465_),
    .A2(_01900_),
    .ZN(_01901_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05320_ (.I0(\u_cpu.rf_ram.memory[132][3] ),
    .I1(\u_cpu.rf_ram.memory[133][3] ),
    .I2(\u_cpu.rf_ram.memory[134][3] ),
    .I3(\u_cpu.rf_ram.memory[135][3] ),
    .S0(_01634_),
    .S1(_01635_),
    .Z(_01902_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05321_ (.A1(_01638_),
    .A2(_01902_),
    .B(_01482_),
    .ZN(_01903_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05322_ (.I0(\u_cpu.rf_ram.memory[136][3] ),
    .I1(\u_cpu.rf_ram.memory[137][3] ),
    .I2(\u_cpu.rf_ram.memory[138][3] ),
    .I3(\u_cpu.rf_ram.memory[139][3] ),
    .S0(_01641_),
    .S1(_01642_),
    .Z(_01904_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05323_ (.A1(_01465_),
    .A2(_01904_),
    .ZN(_01905_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05324_ (.I0(\u_cpu.rf_ram.memory[140][3] ),
    .I1(\u_cpu.rf_ram.memory[141][3] ),
    .I2(\u_cpu.rf_ram.memory[142][3] ),
    .I3(\u_cpu.rf_ram.memory[143][3] ),
    .S0(_01641_),
    .S1(_01642_),
    .Z(_01906_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05325_ (.A1(_01638_),
    .A2(_01906_),
    .B(_01534_),
    .ZN(_01907_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _05326_ (.A1(_01901_),
    .A2(_01903_),
    .B1(_01905_),
    .B2(_01907_),
    .C(_01466_),
    .ZN(_01908_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05327_ (.A1(_01899_),
    .A2(_01908_),
    .ZN(_01909_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05328_ (.A1(_01473_),
    .A2(_01860_),
    .B(_01909_),
    .ZN(_00003_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05329_ (.I0(\u_cpu.rf_ram.memory[28][4] ),
    .I1(\u_cpu.rf_ram.memory[29][4] ),
    .I2(\u_cpu.rf_ram.memory[30][4] ),
    .I3(\u_cpu.rf_ram.memory[31][4] ),
    .S0(_01497_),
    .S1(_01501_),
    .Z(_01910_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05330_ (.A1(_01493_),
    .A2(_01910_),
    .ZN(_01911_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05331_ (.I0(\u_cpu.rf_ram.memory[24][4] ),
    .I1(\u_cpu.rf_ram.memory[25][4] ),
    .I2(\u_cpu.rf_ram.memory[26][4] ),
    .I3(\u_cpu.rf_ram.memory[27][4] ),
    .S0(_01508_),
    .S1(_01509_),
    .Z(_01912_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05332_ (.A1(_01506_),
    .A2(_01912_),
    .B(_01481_),
    .ZN(_01913_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05333_ (.I0(\u_cpu.rf_ram.memory[20][4] ),
    .I1(\u_cpu.rf_ram.memory[21][4] ),
    .I2(\u_cpu.rf_ram.memory[22][4] ),
    .I3(\u_cpu.rf_ram.memory[23][4] ),
    .S0(_01497_),
    .S1(_01501_),
    .Z(_01914_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05334_ (.A1(_01513_),
    .A2(_01914_),
    .ZN(_01915_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05335_ (.I0(\u_cpu.rf_ram.memory[16][4] ),
    .I1(\u_cpu.rf_ram.memory[17][4] ),
    .I2(\u_cpu.rf_ram.memory[18][4] ),
    .I3(\u_cpu.rf_ram.memory[19][4] ),
    .S0(_01508_),
    .S1(_01509_),
    .Z(_01916_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05336_ (.A1(_01506_),
    .A2(_01916_),
    .B(_01519_),
    .ZN(_01917_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _05337_ (.A1(_01911_),
    .A2(_01913_),
    .B1(_01915_),
    .B2(_01917_),
    .C(_01486_),
    .ZN(_01918_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05338_ (.I0(\u_cpu.rf_ram.memory[4][4] ),
    .I1(\u_cpu.rf_ram.memory[5][4] ),
    .I2(\u_cpu.rf_ram.memory[6][4] ),
    .I3(\u_cpu.rf_ram.memory[7][4] ),
    .S0(_01523_),
    .S1(_01525_),
    .Z(_01919_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05339_ (.A1(_01493_),
    .A2(_01919_),
    .ZN(_01920_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05340_ (.I0(\u_cpu.rf_ram.memory[0][4] ),
    .I1(\u_cpu.rf_ram.memory[1][4] ),
    .I2(\u_cpu.rf_ram.memory[2][4] ),
    .I3(\u_cpu.rf_ram.memory[3][4] ),
    .S0(_01530_),
    .S1(_01532_),
    .Z(_01921_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05341_ (.A1(_01528_),
    .A2(_01921_),
    .B(_01534_),
    .ZN(_01922_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05342_ (.I0(\u_cpu.rf_ram.memory[8][4] ),
    .I1(\u_cpu.rf_ram.memory[9][4] ),
    .I2(\u_cpu.rf_ram.memory[10][4] ),
    .I3(\u_cpu.rf_ram.memory[11][4] ),
    .S0(_01523_),
    .S1(_01525_),
    .Z(_01923_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05343_ (.A1(_01528_),
    .A2(_01923_),
    .ZN(_01924_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05344_ (.I0(\u_cpu.rf_ram.memory[12][4] ),
    .I1(\u_cpu.rf_ram.memory[13][4] ),
    .I2(\u_cpu.rf_ram.memory[14][4] ),
    .I3(\u_cpu.rf_ram.memory[15][4] ),
    .S0(_01530_),
    .S1(_01532_),
    .Z(_01925_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05345_ (.A1(_01513_),
    .A2(_01925_),
    .B(_01482_),
    .ZN(_01926_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _05346_ (.A1(_01920_),
    .A2(_01922_),
    .B1(_01924_),
    .B2(_01926_),
    .C(_01541_),
    .ZN(_01927_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05347_ (.I0(\u_cpu.rf_ram.memory[36][4] ),
    .I1(\u_cpu.rf_ram.memory[37][4] ),
    .I2(\u_cpu.rf_ram.memory[38][4] ),
    .I3(\u_cpu.rf_ram.memory[39][4] ),
    .S0(_01544_),
    .S1(_01545_),
    .Z(_01928_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05348_ (.A1(_01543_),
    .A2(_01928_),
    .ZN(_01929_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05349_ (.I0(\u_cpu.rf_ram.memory[32][4] ),
    .I1(\u_cpu.rf_ram.memory[33][4] ),
    .I2(\u_cpu.rf_ram.memory[34][4] ),
    .I3(\u_cpu.rf_ram.memory[35][4] ),
    .S0(_01495_),
    .S1(_01499_),
    .Z(_01930_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05350_ (.A1(_01548_),
    .A2(_01930_),
    .B(_01518_),
    .ZN(_01931_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05351_ (.I0(\u_cpu.rf_ram.memory[40][4] ),
    .I1(\u_cpu.rf_ram.memory[41][4] ),
    .I2(\u_cpu.rf_ram.memory[42][4] ),
    .I3(\u_cpu.rf_ram.memory[43][4] ),
    .S0(_01551_),
    .S1(_01524_),
    .Z(_01932_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05352_ (.A1(_01505_),
    .A2(_01932_),
    .ZN(_01933_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05353_ (.I0(\u_cpu.rf_ram.memory[44][4] ),
    .I1(\u_cpu.rf_ram.memory[45][4] ),
    .I2(\u_cpu.rf_ram.memory[46][4] ),
    .I3(\u_cpu.rf_ram.memory[47][4] ),
    .S0(_01555_),
    .S1(_01531_),
    .Z(_01934_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05354_ (.A1(_01463_),
    .A2(_01934_),
    .B(_01558_),
    .ZN(_01935_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _05355_ (.A1(_01929_),
    .A2(_01931_),
    .B1(_01933_),
    .B2(_01935_),
    .C(_01560_),
    .ZN(_01936_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05356_ (.I0(\u_cpu.rf_ram.memory[60][4] ),
    .I1(\u_cpu.rf_ram.memory[61][4] ),
    .I2(\u_cpu.rf_ram.memory[62][4] ),
    .I3(\u_cpu.rf_ram.memory[63][4] ),
    .S0(_01496_),
    .S1(_01594_),
    .Z(_01937_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05357_ (.A1(_01464_),
    .A2(_01937_),
    .ZN(_01938_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05358_ (.I0(\u_cpu.rf_ram.memory[56][4] ),
    .I1(\u_cpu.rf_ram.memory[57][4] ),
    .I2(\u_cpu.rf_ram.memory[58][4] ),
    .I3(\u_cpu.rf_ram.memory[59][4] ),
    .S0(_01567_),
    .S1(_01568_),
    .Z(_01939_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05359_ (.A1(_01566_),
    .A2(_01939_),
    .B(_01480_),
    .ZN(_01940_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05360_ (.I0(\u_cpu.rf_ram.memory[52][4] ),
    .I1(\u_cpu.rf_ram.memory[53][4] ),
    .I2(\u_cpu.rf_ram.memory[54][4] ),
    .I3(\u_cpu.rf_ram.memory[55][4] ),
    .S0(_01572_),
    .S1(_01573_),
    .Z(_01941_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05361_ (.A1(_01571_),
    .A2(_01941_),
    .ZN(_01942_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05362_ (.I0(\u_cpu.rf_ram.memory[48][4] ),
    .I1(\u_cpu.rf_ram.memory[49][4] ),
    .I2(\u_cpu.rf_ram.memory[50][4] ),
    .I3(\u_cpu.rf_ram.memory[51][4] ),
    .S0(_01576_),
    .S1(_01577_),
    .Z(_01943_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05363_ (.A1(_01505_),
    .A2(_01943_),
    .B(_01579_),
    .ZN(_01944_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _05364_ (.A1(_01938_),
    .A2(_01940_),
    .B1(_01942_),
    .B2(_01944_),
    .C(_01581_),
    .ZN(_01945_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _05365_ (.A1(_01490_),
    .A2(_01936_),
    .A3(_01945_),
    .Z(_01946_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _05366_ (.A1(_01492_),
    .A2(_01918_),
    .A3(_01927_),
    .B(_01946_),
    .ZN(_01947_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05367_ (.I0(\u_cpu.rf_ram.memory[100][4] ),
    .I1(\u_cpu.rf_ram.memory[101][4] ),
    .I2(\u_cpu.rf_ram.memory[102][4] ),
    .I3(\u_cpu.rf_ram.memory[103][4] ),
    .S0(_01551_),
    .S1(_01524_),
    .Z(_01948_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05368_ (.A1(_01571_),
    .A2(_01948_),
    .ZN(_01949_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05369_ (.I0(\u_cpu.rf_ram.memory[96][4] ),
    .I1(\u_cpu.rf_ram.memory[97][4] ),
    .I2(\u_cpu.rf_ram.memory[98][4] ),
    .I3(\u_cpu.rf_ram.memory[99][4] ),
    .S0(_01567_),
    .S1(_01568_),
    .Z(_01950_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05370_ (.A1(_01548_),
    .A2(_01950_),
    .B(_01579_),
    .ZN(_01951_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05371_ (.I0(\u_cpu.rf_ram.memory[108][4] ),
    .I1(\u_cpu.rf_ram.memory[109][4] ),
    .I2(\u_cpu.rf_ram.memory[110][4] ),
    .I3(\u_cpu.rf_ram.memory[111][4] ),
    .S0(_01529_),
    .S1(_01500_),
    .Z(_01952_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05372_ (.A1(_01512_),
    .A2(_01952_),
    .ZN(_01953_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05373_ (.I0(\u_cpu.rf_ram.memory[104][4] ),
    .I1(\u_cpu.rf_ram.memory[105][4] ),
    .I2(\u_cpu.rf_ram.memory[106][4] ),
    .I3(\u_cpu.rf_ram.memory[107][4] ),
    .S0(_01555_),
    .S1(_01531_),
    .Z(_01954_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05374_ (.A1(_01566_),
    .A2(_01954_),
    .B(_01558_),
    .ZN(_01955_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _05375_ (.A1(_01949_),
    .A2(_01951_),
    .B1(_01953_),
    .B2(_01955_),
    .C(_01560_),
    .ZN(_01956_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05376_ (.I0(\u_cpu.rf_ram.memory[124][4] ),
    .I1(\u_cpu.rf_ram.memory[125][4] ),
    .I2(\u_cpu.rf_ram.memory[126][4] ),
    .I3(\u_cpu.rf_ram.memory[127][4] ),
    .S0(_01496_),
    .S1(_01594_),
    .Z(_01957_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05377_ (.A1(_01543_),
    .A2(_01957_),
    .ZN(_01958_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05378_ (.I0(\u_cpu.rf_ram.memory[120][4] ),
    .I1(\u_cpu.rf_ram.memory[121][4] ),
    .I2(\u_cpu.rf_ram.memory[122][4] ),
    .I3(\u_cpu.rf_ram.memory[123][4] ),
    .S0(_01598_),
    .S1(_01556_),
    .Z(_01959_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05379_ (.A1(_01597_),
    .A2(_01959_),
    .B(_01600_),
    .ZN(_01960_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05380_ (.I0(\u_cpu.rf_ram.memory[112][4] ),
    .I1(\u_cpu.rf_ram.memory[113][4] ),
    .I2(\u_cpu.rf_ram.memory[114][4] ),
    .I3(\u_cpu.rf_ram.memory[115][4] ),
    .S0(_01572_),
    .S1(_01573_),
    .Z(_01961_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05381_ (.A1(_01602_),
    .A2(_01961_),
    .ZN(_01962_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05382_ (.I0(\u_cpu.rf_ram.memory[116][4] ),
    .I1(\u_cpu.rf_ram.memory[117][4] ),
    .I2(\u_cpu.rf_ram.memory[118][4] ),
    .I3(\u_cpu.rf_ram.memory[119][4] ),
    .S0(_01576_),
    .S1(_01577_),
    .Z(_01963_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05383_ (.A1(_01554_),
    .A2(_01963_),
    .B(_01607_),
    .ZN(_01964_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _05384_ (.A1(_01958_),
    .A2(_01960_),
    .B1(_01962_),
    .B2(_01964_),
    .C(_01581_),
    .ZN(_01965_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _05385_ (.A1(_01490_),
    .A2(_01956_),
    .A3(_01965_),
    .ZN(_01966_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05386_ (.I0(\u_cpu.rf_ram.memory[92][4] ),
    .I1(\u_cpu.rf_ram.memory[93][4] ),
    .I2(\u_cpu.rf_ram.memory[94][4] ),
    .I3(\u_cpu.rf_ram.memory[95][4] ),
    .S0(_01562_),
    .S1(_01563_),
    .Z(_01967_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05387_ (.A1(_01464_),
    .A2(_01967_),
    .ZN(_01968_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05388_ (.I0(\u_cpu.rf_ram.memory[88][4] ),
    .I1(\u_cpu.rf_ram.memory[89][4] ),
    .I2(\u_cpu.rf_ram.memory[90][4] ),
    .I3(\u_cpu.rf_ram.memory[91][4] ),
    .S0(_01598_),
    .S1(_01556_),
    .Z(_01969_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05389_ (.A1(_01597_),
    .A2(_01969_),
    .B(_01600_),
    .ZN(_01970_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05390_ (.I0(\u_cpu.rf_ram.memory[80][4] ),
    .I1(\u_cpu.rf_ram.memory[81][4] ),
    .I2(\u_cpu.rf_ram.memory[82][4] ),
    .I3(\u_cpu.rf_ram.memory[83][4] ),
    .S0(_01544_),
    .S1(_01545_),
    .Z(_01971_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05391_ (.A1(_01602_),
    .A2(_01971_),
    .ZN(_01972_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05392_ (.I0(\u_cpu.rf_ram.memory[84][4] ),
    .I1(\u_cpu.rf_ram.memory[85][4] ),
    .I2(\u_cpu.rf_ram.memory[86][4] ),
    .I3(\u_cpu.rf_ram.memory[87][4] ),
    .S0(_01507_),
    .S1(_01605_),
    .Z(_01973_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05393_ (.A1(_01554_),
    .A2(_01973_),
    .B(_01607_),
    .ZN(_01974_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _05394_ (.A1(_01968_),
    .A2(_01970_),
    .B1(_01972_),
    .B2(_01974_),
    .C(_01486_),
    .ZN(_01975_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05395_ (.I0(\u_cpu.rf_ram.memory[64][4] ),
    .I1(\u_cpu.rf_ram.memory[65][4] ),
    .I2(\u_cpu.rf_ram.memory[66][4] ),
    .I3(\u_cpu.rf_ram.memory[67][4] ),
    .S0(_01522_),
    .S1(_01622_),
    .Z(_01976_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05396_ (.A1(_01621_),
    .A2(_01976_),
    .ZN(_01977_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05397_ (.I0(\u_cpu.rf_ram.memory[68][4] ),
    .I1(\u_cpu.rf_ram.memory[69][4] ),
    .I2(\u_cpu.rf_ram.memory[70][4] ),
    .I3(\u_cpu.rf_ram.memory[71][4] ),
    .S0(_01507_),
    .S1(_01605_),
    .Z(_01978_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05398_ (.A1(_01617_),
    .A2(_01978_),
    .B(_01519_),
    .ZN(_01979_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05399_ (.I0(\u_cpu.rf_ram.memory[72][4] ),
    .I1(\u_cpu.rf_ram.memory[73][4] ),
    .I2(\u_cpu.rf_ram.memory[74][4] ),
    .I3(\u_cpu.rf_ram.memory[75][4] ),
    .S0(_01562_),
    .S1(_01622_),
    .Z(_01980_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05400_ (.A1(_01621_),
    .A2(_01980_),
    .ZN(_01981_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05401_ (.I0(\u_cpu.rf_ram.memory[76][4] ),
    .I1(\u_cpu.rf_ram.memory[77][4] ),
    .I2(\u_cpu.rf_ram.memory[78][4] ),
    .I3(\u_cpu.rf_ram.memory[79][4] ),
    .S0(_01529_),
    .S1(_01500_),
    .Z(_01982_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05402_ (.A1(_01617_),
    .A2(_01982_),
    .B(_01481_),
    .ZN(_01983_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _05403_ (.A1(_01977_),
    .A2(_01979_),
    .B1(_01981_),
    .B2(_01983_),
    .C(_01541_),
    .ZN(_01984_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _05404_ (.A1(_01492_),
    .A2(_01975_),
    .A3(_01984_),
    .ZN(_01985_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05405_ (.A1(_01966_),
    .A2(_01985_),
    .B(_01471_),
    .ZN(_01986_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05406_ (.I0(\u_cpu.rf_ram.memory[136][4] ),
    .I1(\u_cpu.rf_ram.memory[137][4] ),
    .I2(\u_cpu.rf_ram.memory[138][4] ),
    .I3(\u_cpu.rf_ram.memory[139][4] ),
    .S0(_01634_),
    .S1(_01635_),
    .Z(_01987_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05407_ (.A1(_01465_),
    .A2(_01987_),
    .ZN(_01988_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05408_ (.I0(\u_cpu.rf_ram.memory[140][4] ),
    .I1(\u_cpu.rf_ram.memory[141][4] ),
    .I2(\u_cpu.rf_ram.memory[142][4] ),
    .I3(\u_cpu.rf_ram.memory[143][4] ),
    .S0(_01634_),
    .S1(_01635_),
    .Z(_01989_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05409_ (.A1(_01638_),
    .A2(_01989_),
    .B(_01534_),
    .ZN(_01990_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05410_ (.I0(\u_cpu.rf_ram.memory[128][4] ),
    .I1(\u_cpu.rf_ram.memory[129][4] ),
    .I2(\u_cpu.rf_ram.memory[130][4] ),
    .I3(\u_cpu.rf_ram.memory[131][4] ),
    .S0(_01641_),
    .S1(_01642_),
    .Z(_01991_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05411_ (.A1(_01465_),
    .A2(_01991_),
    .ZN(_01992_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05412_ (.I0(\u_cpu.rf_ram.memory[132][4] ),
    .I1(\u_cpu.rf_ram.memory[133][4] ),
    .I2(\u_cpu.rf_ram.memory[134][4] ),
    .I3(\u_cpu.rf_ram.memory[135][4] ),
    .S0(_01641_),
    .S1(_01642_),
    .Z(_01993_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05413_ (.A1(_01638_),
    .A2(_01993_),
    .B(_01482_),
    .ZN(_01994_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _05414_ (.A1(_01988_),
    .A2(_01990_),
    .B1(_01992_),
    .B2(_01994_),
    .C(_01466_),
    .ZN(_01995_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05415_ (.A1(_01986_),
    .A2(_01995_),
    .ZN(_01996_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05416_ (.A1(_01473_),
    .A2(_01947_),
    .B(_01996_),
    .ZN(_00004_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05417_ (.I0(\u_cpu.rf_ram.memory[28][5] ),
    .I1(\u_cpu.rf_ram.memory[29][5] ),
    .I2(\u_cpu.rf_ram.memory[30][5] ),
    .I3(\u_cpu.rf_ram.memory[31][5] ),
    .S0(_01497_),
    .S1(_01501_),
    .Z(_01997_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05418_ (.A1(_01493_),
    .A2(_01997_),
    .ZN(_01998_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05419_ (.I0(\u_cpu.rf_ram.memory[24][5] ),
    .I1(\u_cpu.rf_ram.memory[25][5] ),
    .I2(\u_cpu.rf_ram.memory[26][5] ),
    .I3(\u_cpu.rf_ram.memory[27][5] ),
    .S0(_01508_),
    .S1(_01509_),
    .Z(_01999_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05420_ (.A1(_01506_),
    .A2(_01999_),
    .B(_01481_),
    .ZN(_02000_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05421_ (.I0(\u_cpu.rf_ram.memory[20][5] ),
    .I1(\u_cpu.rf_ram.memory[21][5] ),
    .I2(\u_cpu.rf_ram.memory[22][5] ),
    .I3(\u_cpu.rf_ram.memory[23][5] ),
    .S0(_01497_),
    .S1(_01501_),
    .Z(_02001_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05422_ (.A1(_01513_),
    .A2(_02001_),
    .ZN(_02002_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05423_ (.I0(\u_cpu.rf_ram.memory[16][5] ),
    .I1(\u_cpu.rf_ram.memory[17][5] ),
    .I2(\u_cpu.rf_ram.memory[18][5] ),
    .I3(\u_cpu.rf_ram.memory[19][5] ),
    .S0(_01508_),
    .S1(_01509_),
    .Z(_02003_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05424_ (.A1(_01506_),
    .A2(_02003_),
    .B(_01519_),
    .ZN(_02004_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _05425_ (.A1(_01998_),
    .A2(_02000_),
    .B1(_02002_),
    .B2(_02004_),
    .C(_01486_),
    .ZN(_02005_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05426_ (.I0(\u_cpu.rf_ram.memory[4][5] ),
    .I1(\u_cpu.rf_ram.memory[5][5] ),
    .I2(\u_cpu.rf_ram.memory[6][5] ),
    .I3(\u_cpu.rf_ram.memory[7][5] ),
    .S0(_01523_),
    .S1(_01525_),
    .Z(_02006_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05427_ (.A1(_01493_),
    .A2(_02006_),
    .ZN(_02007_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05428_ (.I0(\u_cpu.rf_ram.memory[0][5] ),
    .I1(\u_cpu.rf_ram.memory[1][5] ),
    .I2(\u_cpu.rf_ram.memory[2][5] ),
    .I3(\u_cpu.rf_ram.memory[3][5] ),
    .S0(_01530_),
    .S1(_01532_),
    .Z(_02008_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05429_ (.A1(_01528_),
    .A2(_02008_),
    .B(_01534_),
    .ZN(_02009_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05430_ (.I0(\u_cpu.rf_ram.memory[8][5] ),
    .I1(\u_cpu.rf_ram.memory[9][5] ),
    .I2(\u_cpu.rf_ram.memory[10][5] ),
    .I3(\u_cpu.rf_ram.memory[11][5] ),
    .S0(_01523_),
    .S1(_01525_),
    .Z(_02010_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05431_ (.A1(_01528_),
    .A2(_02010_),
    .ZN(_02011_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05432_ (.I0(\u_cpu.rf_ram.memory[12][5] ),
    .I1(\u_cpu.rf_ram.memory[13][5] ),
    .I2(\u_cpu.rf_ram.memory[14][5] ),
    .I3(\u_cpu.rf_ram.memory[15][5] ),
    .S0(_01530_),
    .S1(_01532_),
    .Z(_02012_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05433_ (.A1(_01513_),
    .A2(_02012_),
    .B(_01482_),
    .ZN(_02013_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _05434_ (.A1(_02007_),
    .A2(_02009_),
    .B1(_02011_),
    .B2(_02013_),
    .C(_01541_),
    .ZN(_02014_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05435_ (.I0(\u_cpu.rf_ram.memory[36][5] ),
    .I1(\u_cpu.rf_ram.memory[37][5] ),
    .I2(\u_cpu.rf_ram.memory[38][5] ),
    .I3(\u_cpu.rf_ram.memory[39][5] ),
    .S0(_01544_),
    .S1(_01545_),
    .Z(_02015_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05436_ (.A1(_01571_),
    .A2(_02015_),
    .ZN(_02016_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05437_ (.I0(\u_cpu.rf_ram.memory[32][5] ),
    .I1(\u_cpu.rf_ram.memory[33][5] ),
    .I2(\u_cpu.rf_ram.memory[34][5] ),
    .I3(\u_cpu.rf_ram.memory[35][5] ),
    .S0(_01495_),
    .S1(_01499_),
    .Z(_02017_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05438_ (.A1(_01504_),
    .A2(_02017_),
    .B(_01518_),
    .ZN(_02018_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05439_ (.I0(\u_cpu.rf_ram.memory[40][5] ),
    .I1(\u_cpu.rf_ram.memory[41][5] ),
    .I2(\u_cpu.rf_ram.memory[42][5] ),
    .I3(\u_cpu.rf_ram.memory[43][5] ),
    .S0(_01551_),
    .S1(_01524_),
    .Z(_02019_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05440_ (.A1(_01505_),
    .A2(_02019_),
    .ZN(_02020_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05441_ (.I0(\u_cpu.rf_ram.memory[44][5] ),
    .I1(\u_cpu.rf_ram.memory[45][5] ),
    .I2(\u_cpu.rf_ram.memory[46][5] ),
    .I3(\u_cpu.rf_ram.memory[47][5] ),
    .S0(_01555_),
    .S1(_01531_),
    .Z(_02021_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05442_ (.A1(_01463_),
    .A2(_02021_),
    .B(_01558_),
    .ZN(_02022_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _05443_ (.A1(_02016_),
    .A2(_02018_),
    .B1(_02020_),
    .B2(_02022_),
    .C(_01560_),
    .ZN(_02023_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05444_ (.I0(\u_cpu.rf_ram.memory[60][5] ),
    .I1(\u_cpu.rf_ram.memory[61][5] ),
    .I2(\u_cpu.rf_ram.memory[62][5] ),
    .I3(\u_cpu.rf_ram.memory[63][5] ),
    .S0(_01496_),
    .S1(_01594_),
    .Z(_02024_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05445_ (.A1(_01543_),
    .A2(_02024_),
    .ZN(_02025_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05446_ (.I0(\u_cpu.rf_ram.memory[56][5] ),
    .I1(\u_cpu.rf_ram.memory[57][5] ),
    .I2(\u_cpu.rf_ram.memory[58][5] ),
    .I3(\u_cpu.rf_ram.memory[59][5] ),
    .S0(_01567_),
    .S1(_01568_),
    .Z(_02026_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05447_ (.A1(_01548_),
    .A2(_02026_),
    .B(_01480_),
    .ZN(_02027_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05448_ (.I0(\u_cpu.rf_ram.memory[52][5] ),
    .I1(\u_cpu.rf_ram.memory[53][5] ),
    .I2(\u_cpu.rf_ram.memory[54][5] ),
    .I3(\u_cpu.rf_ram.memory[55][5] ),
    .S0(_01572_),
    .S1(_01573_),
    .Z(_02028_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05449_ (.A1(_01571_),
    .A2(_02028_),
    .ZN(_02029_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05450_ (.I0(\u_cpu.rf_ram.memory[48][5] ),
    .I1(\u_cpu.rf_ram.memory[49][5] ),
    .I2(\u_cpu.rf_ram.memory[50][5] ),
    .I3(\u_cpu.rf_ram.memory[51][5] ),
    .S0(_01576_),
    .S1(_01577_),
    .Z(_02030_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05451_ (.A1(_01597_),
    .A2(_02030_),
    .B(_01579_),
    .ZN(_02031_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _05452_ (.A1(_02025_),
    .A2(_02027_),
    .B1(_02029_),
    .B2(_02031_),
    .C(_01581_),
    .ZN(_02032_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _05453_ (.A1(_01490_),
    .A2(_02023_),
    .A3(_02032_),
    .Z(_02033_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _05454_ (.A1(_01492_),
    .A2(_02005_),
    .A3(_02014_),
    .B(_02033_),
    .ZN(_02034_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05455_ (.I0(\u_cpu.rf_ram.memory[100][5] ),
    .I1(\u_cpu.rf_ram.memory[101][5] ),
    .I2(\u_cpu.rf_ram.memory[102][5] ),
    .I3(\u_cpu.rf_ram.memory[103][5] ),
    .S0(_01551_),
    .S1(_01524_),
    .Z(_02035_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05456_ (.A1(_01512_),
    .A2(_02035_),
    .ZN(_02036_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05457_ (.I0(\u_cpu.rf_ram.memory[96][5] ),
    .I1(\u_cpu.rf_ram.memory[97][5] ),
    .I2(\u_cpu.rf_ram.memory[98][5] ),
    .I3(\u_cpu.rf_ram.memory[99][5] ),
    .S0(_01567_),
    .S1(_01568_),
    .Z(_02037_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05458_ (.A1(_01548_),
    .A2(_02037_),
    .B(_01579_),
    .ZN(_02038_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05459_ (.I0(\u_cpu.rf_ram.memory[108][5] ),
    .I1(\u_cpu.rf_ram.memory[109][5] ),
    .I2(\u_cpu.rf_ram.memory[110][5] ),
    .I3(\u_cpu.rf_ram.memory[111][5] ),
    .S0(_01529_),
    .S1(_01500_),
    .Z(_02039_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05460_ (.A1(_01512_),
    .A2(_02039_),
    .ZN(_02040_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05461_ (.I0(\u_cpu.rf_ram.memory[104][5] ),
    .I1(\u_cpu.rf_ram.memory[105][5] ),
    .I2(\u_cpu.rf_ram.memory[106][5] ),
    .I3(\u_cpu.rf_ram.memory[107][5] ),
    .S0(_01555_),
    .S1(_01531_),
    .Z(_02041_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05462_ (.A1(_01566_),
    .A2(_02041_),
    .B(_01558_),
    .ZN(_02042_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _05463_ (.A1(_02036_),
    .A2(_02038_),
    .B1(_02040_),
    .B2(_02042_),
    .C(_01560_),
    .ZN(_02043_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05464_ (.I0(\u_cpu.rf_ram.memory[124][5] ),
    .I1(\u_cpu.rf_ram.memory[125][5] ),
    .I2(\u_cpu.rf_ram.memory[126][5] ),
    .I3(\u_cpu.rf_ram.memory[127][5] ),
    .S0(_01496_),
    .S1(_01594_),
    .Z(_02044_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05465_ (.A1(_01543_),
    .A2(_02044_),
    .ZN(_02045_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05466_ (.I0(\u_cpu.rf_ram.memory[120][5] ),
    .I1(\u_cpu.rf_ram.memory[121][5] ),
    .I2(\u_cpu.rf_ram.memory[122][5] ),
    .I3(\u_cpu.rf_ram.memory[123][5] ),
    .S0(_01598_),
    .S1(_01556_),
    .Z(_02046_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05467_ (.A1(_01566_),
    .A2(_02046_),
    .B(_01600_),
    .ZN(_02047_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05468_ (.I0(\u_cpu.rf_ram.memory[112][5] ),
    .I1(\u_cpu.rf_ram.memory[113][5] ),
    .I2(\u_cpu.rf_ram.memory[114][5] ),
    .I3(\u_cpu.rf_ram.memory[115][5] ),
    .S0(_01572_),
    .S1(_01573_),
    .Z(_02048_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05469_ (.A1(_01602_),
    .A2(_02048_),
    .ZN(_02049_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05470_ (.I0(\u_cpu.rf_ram.memory[116][5] ),
    .I1(\u_cpu.rf_ram.memory[117][5] ),
    .I2(\u_cpu.rf_ram.memory[118][5] ),
    .I3(\u_cpu.rf_ram.memory[119][5] ),
    .S0(_01576_),
    .S1(_01577_),
    .Z(_02050_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05471_ (.A1(_01554_),
    .A2(_02050_),
    .B(_01607_),
    .ZN(_02051_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _05472_ (.A1(_02045_),
    .A2(_02047_),
    .B1(_02049_),
    .B2(_02051_),
    .C(_01581_),
    .ZN(_02052_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _05473_ (.A1(_01490_),
    .A2(_02043_),
    .A3(_02052_),
    .ZN(_02053_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05474_ (.I0(\u_cpu.rf_ram.memory[92][5] ),
    .I1(\u_cpu.rf_ram.memory[93][5] ),
    .I2(\u_cpu.rf_ram.memory[94][5] ),
    .I3(\u_cpu.rf_ram.memory[95][5] ),
    .S0(_01562_),
    .S1(_01563_),
    .Z(_02054_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05475_ (.A1(_01464_),
    .A2(_02054_),
    .ZN(_02055_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05476_ (.I0(\u_cpu.rf_ram.memory[88][5] ),
    .I1(\u_cpu.rf_ram.memory[89][5] ),
    .I2(\u_cpu.rf_ram.memory[90][5] ),
    .I3(\u_cpu.rf_ram.memory[91][5] ),
    .S0(_01598_),
    .S1(_01556_),
    .Z(_02056_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05477_ (.A1(_01597_),
    .A2(_02056_),
    .B(_01600_),
    .ZN(_02057_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05478_ (.I0(\u_cpu.rf_ram.memory[80][5] ),
    .I1(\u_cpu.rf_ram.memory[81][5] ),
    .I2(\u_cpu.rf_ram.memory[82][5] ),
    .I3(\u_cpu.rf_ram.memory[83][5] ),
    .S0(_01544_),
    .S1(_01545_),
    .Z(_02058_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05479_ (.A1(_01602_),
    .A2(_02058_),
    .ZN(_02059_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05480_ (.I0(\u_cpu.rf_ram.memory[84][5] ),
    .I1(\u_cpu.rf_ram.memory[85][5] ),
    .I2(\u_cpu.rf_ram.memory[86][5] ),
    .I3(\u_cpu.rf_ram.memory[87][5] ),
    .S0(_01507_),
    .S1(_01605_),
    .Z(_02060_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05481_ (.A1(_01554_),
    .A2(_02060_),
    .B(_01607_),
    .ZN(_02061_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _05482_ (.A1(_02055_),
    .A2(_02057_),
    .B1(_02059_),
    .B2(_02061_),
    .C(_01486_),
    .ZN(_02062_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05483_ (.I0(\u_cpu.rf_ram.memory[64][5] ),
    .I1(\u_cpu.rf_ram.memory[65][5] ),
    .I2(\u_cpu.rf_ram.memory[66][5] ),
    .I3(\u_cpu.rf_ram.memory[67][5] ),
    .S0(_01522_),
    .S1(_01622_),
    .Z(_02063_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05484_ (.A1(_01621_),
    .A2(_02063_),
    .ZN(_02064_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05485_ (.I0(\u_cpu.rf_ram.memory[68][5] ),
    .I1(\u_cpu.rf_ram.memory[69][5] ),
    .I2(\u_cpu.rf_ram.memory[70][5] ),
    .I3(\u_cpu.rf_ram.memory[71][5] ),
    .S0(_01507_),
    .S1(_01605_),
    .Z(_02065_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05486_ (.A1(_01617_),
    .A2(_02065_),
    .B(_01519_),
    .ZN(_02066_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05487_ (.I0(\u_cpu.rf_ram.memory[72][5] ),
    .I1(\u_cpu.rf_ram.memory[73][5] ),
    .I2(\u_cpu.rf_ram.memory[74][5] ),
    .I3(\u_cpu.rf_ram.memory[75][5] ),
    .S0(_01562_),
    .S1(_01563_),
    .Z(_02067_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05488_ (.A1(_01621_),
    .A2(_02067_),
    .ZN(_02068_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05489_ (.I0(\u_cpu.rf_ram.memory[76][5] ),
    .I1(\u_cpu.rf_ram.memory[77][5] ),
    .I2(\u_cpu.rf_ram.memory[78][5] ),
    .I3(\u_cpu.rf_ram.memory[79][5] ),
    .S0(_01529_),
    .S1(_01500_),
    .Z(_02069_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05490_ (.A1(_01617_),
    .A2(_02069_),
    .B(_01481_),
    .ZN(_02070_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _05491_ (.A1(_02064_),
    .A2(_02066_),
    .B1(_02068_),
    .B2(_02070_),
    .C(_01541_),
    .ZN(_02071_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _05492_ (.A1(_01492_),
    .A2(_02062_),
    .A3(_02071_),
    .ZN(_02072_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05493_ (.A1(_02053_),
    .A2(_02072_),
    .B(_01471_),
    .ZN(_02073_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05494_ (.I0(\u_cpu.rf_ram.memory[136][5] ),
    .I1(\u_cpu.rf_ram.memory[137][5] ),
    .I2(\u_cpu.rf_ram.memory[138][5] ),
    .I3(\u_cpu.rf_ram.memory[139][5] ),
    .S0(_01634_),
    .S1(_01635_),
    .Z(_02074_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05495_ (.A1(_01465_),
    .A2(_02074_),
    .ZN(_02075_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05496_ (.I0(\u_cpu.rf_ram.memory[140][5] ),
    .I1(\u_cpu.rf_ram.memory[141][5] ),
    .I2(\u_cpu.rf_ram.memory[142][5] ),
    .I3(\u_cpu.rf_ram.memory[143][5] ),
    .S0(_01634_),
    .S1(_01635_),
    .Z(_02076_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05497_ (.A1(_01638_),
    .A2(_02076_),
    .B(_01534_),
    .ZN(_02077_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05498_ (.I0(\u_cpu.rf_ram.memory[128][5] ),
    .I1(\u_cpu.rf_ram.memory[129][5] ),
    .I2(\u_cpu.rf_ram.memory[130][5] ),
    .I3(\u_cpu.rf_ram.memory[131][5] ),
    .S0(_01641_),
    .S1(_01642_),
    .Z(_02078_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05499_ (.A1(_01465_),
    .A2(_02078_),
    .ZN(_02079_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05500_ (.I0(\u_cpu.rf_ram.memory[132][5] ),
    .I1(\u_cpu.rf_ram.memory[133][5] ),
    .I2(\u_cpu.rf_ram.memory[134][5] ),
    .I3(\u_cpu.rf_ram.memory[135][5] ),
    .S0(_01641_),
    .S1(_01642_),
    .Z(_02080_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05501_ (.A1(_01638_),
    .A2(_02080_),
    .B(_01482_),
    .ZN(_02081_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _05502_ (.A1(_02075_),
    .A2(_02077_),
    .B1(_02079_),
    .B2(_02081_),
    .C(_01466_),
    .ZN(_02082_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05503_ (.A1(_02073_),
    .A2(_02082_),
    .ZN(_02083_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05504_ (.A1(_01473_),
    .A2(_02034_),
    .B(_02083_),
    .ZN(_00005_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05505_ (.I0(\u_cpu.rf_ram.memory[28][6] ),
    .I1(\u_cpu.rf_ram.memory[29][6] ),
    .I2(\u_cpu.rf_ram.memory[30][6] ),
    .I3(\u_cpu.rf_ram.memory[31][6] ),
    .S0(_01497_),
    .S1(_01501_),
    .Z(_02084_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05506_ (.A1(_01493_),
    .A2(_02084_),
    .ZN(_02085_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05507_ (.I0(\u_cpu.rf_ram.memory[24][6] ),
    .I1(\u_cpu.rf_ram.memory[25][6] ),
    .I2(\u_cpu.rf_ram.memory[26][6] ),
    .I3(\u_cpu.rf_ram.memory[27][6] ),
    .S0(_01522_),
    .S1(_01509_),
    .Z(_02086_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05508_ (.A1(_01506_),
    .A2(_02086_),
    .B(_01481_),
    .ZN(_02087_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05509_ (.I0(\u_cpu.rf_ram.memory[20][6] ),
    .I1(\u_cpu.rf_ram.memory[21][6] ),
    .I2(\u_cpu.rf_ram.memory[22][6] ),
    .I3(\u_cpu.rf_ram.memory[23][6] ),
    .S0(_01530_),
    .S1(_01501_),
    .Z(_02088_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05510_ (.A1(_01513_),
    .A2(_02088_),
    .ZN(_02089_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05511_ (.I0(\u_cpu.rf_ram.memory[16][6] ),
    .I1(\u_cpu.rf_ram.memory[17][6] ),
    .I2(\u_cpu.rf_ram.memory[18][6] ),
    .I3(\u_cpu.rf_ram.memory[19][6] ),
    .S0(_01508_),
    .S1(_01509_),
    .Z(_02090_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05512_ (.A1(_01506_),
    .A2(_02090_),
    .B(_01519_),
    .ZN(_02091_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _05513_ (.A1(_02085_),
    .A2(_02087_),
    .B1(_02089_),
    .B2(_02091_),
    .C(_01486_),
    .ZN(_02092_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05514_ (.I0(\u_cpu.rf_ram.memory[4][6] ),
    .I1(\u_cpu.rf_ram.memory[5][6] ),
    .I2(\u_cpu.rf_ram.memory[6][6] ),
    .I3(\u_cpu.rf_ram.memory[7][6] ),
    .S0(_01523_),
    .S1(_01525_),
    .Z(_02093_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05515_ (.A1(_01493_),
    .A2(_02093_),
    .ZN(_02094_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05516_ (.I0(\u_cpu.rf_ram.memory[0][6] ),
    .I1(\u_cpu.rf_ram.memory[1][6] ),
    .I2(\u_cpu.rf_ram.memory[2][6] ),
    .I3(\u_cpu.rf_ram.memory[3][6] ),
    .S0(_01508_),
    .S1(_01532_),
    .Z(_02095_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05517_ (.A1(_01528_),
    .A2(_02095_),
    .B(_01534_),
    .ZN(_02096_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05518_ (.I0(\u_cpu.rf_ram.memory[8][6] ),
    .I1(\u_cpu.rf_ram.memory[9][6] ),
    .I2(\u_cpu.rf_ram.memory[10][6] ),
    .I3(\u_cpu.rf_ram.memory[11][6] ),
    .S0(_01497_),
    .S1(_01525_),
    .Z(_02097_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05519_ (.A1(_01528_),
    .A2(_02097_),
    .ZN(_02098_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05520_ (.I0(\u_cpu.rf_ram.memory[12][6] ),
    .I1(\u_cpu.rf_ram.memory[13][6] ),
    .I2(\u_cpu.rf_ram.memory[14][6] ),
    .I3(\u_cpu.rf_ram.memory[15][6] ),
    .S0(_01530_),
    .S1(_01532_),
    .Z(_02099_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05521_ (.A1(_01513_),
    .A2(_02099_),
    .B(_01482_),
    .ZN(_02100_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _05522_ (.A1(_02094_),
    .A2(_02096_),
    .B1(_02098_),
    .B2(_02100_),
    .C(_01541_),
    .ZN(_02101_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05523_ (.I0(\u_cpu.rf_ram.memory[36][6] ),
    .I1(\u_cpu.rf_ram.memory[37][6] ),
    .I2(\u_cpu.rf_ram.memory[38][6] ),
    .I3(\u_cpu.rf_ram.memory[39][6] ),
    .S0(_01544_),
    .S1(_01545_),
    .Z(_02102_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05524_ (.A1(_01571_),
    .A2(_02102_),
    .ZN(_02103_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05525_ (.I0(\u_cpu.rf_ram.memory[32][6] ),
    .I1(\u_cpu.rf_ram.memory[33][6] ),
    .I2(\u_cpu.rf_ram.memory[34][6] ),
    .I3(\u_cpu.rf_ram.memory[35][6] ),
    .S0(_01495_),
    .S1(_01499_),
    .Z(_02104_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05526_ (.A1(_01504_),
    .A2(_02104_),
    .B(_01518_),
    .ZN(_02105_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05527_ (.I0(\u_cpu.rf_ram.memory[40][6] ),
    .I1(\u_cpu.rf_ram.memory[41][6] ),
    .I2(\u_cpu.rf_ram.memory[42][6] ),
    .I3(\u_cpu.rf_ram.memory[43][6] ),
    .S0(_01551_),
    .S1(_01524_),
    .Z(_02106_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05528_ (.A1(_01505_),
    .A2(_02106_),
    .ZN(_02107_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05529_ (.I0(\u_cpu.rf_ram.memory[44][6] ),
    .I1(\u_cpu.rf_ram.memory[45][6] ),
    .I2(\u_cpu.rf_ram.memory[46][6] ),
    .I3(\u_cpu.rf_ram.memory[47][6] ),
    .S0(_01555_),
    .S1(_01531_),
    .Z(_02108_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05530_ (.A1(_01463_),
    .A2(_02108_),
    .B(_01558_),
    .ZN(_02109_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _05531_ (.A1(_02103_),
    .A2(_02105_),
    .B1(_02107_),
    .B2(_02109_),
    .C(_01560_),
    .ZN(_02110_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05532_ (.I0(\u_cpu.rf_ram.memory[60][6] ),
    .I1(\u_cpu.rf_ram.memory[61][6] ),
    .I2(\u_cpu.rf_ram.memory[62][6] ),
    .I3(\u_cpu.rf_ram.memory[63][6] ),
    .S0(_01496_),
    .S1(_01594_),
    .Z(_02111_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05533_ (.A1(_01543_),
    .A2(_02111_),
    .ZN(_02112_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05534_ (.I0(\u_cpu.rf_ram.memory[56][6] ),
    .I1(\u_cpu.rf_ram.memory[57][6] ),
    .I2(\u_cpu.rf_ram.memory[58][6] ),
    .I3(\u_cpu.rf_ram.memory[59][6] ),
    .S0(_01567_),
    .S1(_01568_),
    .Z(_02113_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05535_ (.A1(_01548_),
    .A2(_02113_),
    .B(_01480_),
    .ZN(_02114_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05536_ (.I0(\u_cpu.rf_ram.memory[52][6] ),
    .I1(\u_cpu.rf_ram.memory[53][6] ),
    .I2(\u_cpu.rf_ram.memory[54][6] ),
    .I3(\u_cpu.rf_ram.memory[55][6] ),
    .S0(_01572_),
    .S1(_01573_),
    .Z(_02115_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05537_ (.A1(_01571_),
    .A2(_02115_),
    .ZN(_02116_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05538_ (.I0(\u_cpu.rf_ram.memory[48][6] ),
    .I1(\u_cpu.rf_ram.memory[49][6] ),
    .I2(\u_cpu.rf_ram.memory[50][6] ),
    .I3(\u_cpu.rf_ram.memory[51][6] ),
    .S0(_01576_),
    .S1(_01577_),
    .Z(_02117_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05539_ (.A1(_01597_),
    .A2(_02117_),
    .B(_01579_),
    .ZN(_02118_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _05540_ (.A1(_02112_),
    .A2(_02114_),
    .B1(_02116_),
    .B2(_02118_),
    .C(_01581_),
    .ZN(_02119_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _05541_ (.A1(_01490_),
    .A2(_02110_),
    .A3(_02119_),
    .Z(_02120_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _05542_ (.A1(_01492_),
    .A2(_02092_),
    .A3(_02101_),
    .B(_02120_),
    .ZN(_02121_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05543_ (.I0(\u_cpu.rf_ram.memory[100][6] ),
    .I1(\u_cpu.rf_ram.memory[101][6] ),
    .I2(\u_cpu.rf_ram.memory[102][6] ),
    .I3(\u_cpu.rf_ram.memory[103][6] ),
    .S0(_01551_),
    .S1(_01524_),
    .Z(_02122_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05544_ (.A1(_01512_),
    .A2(_02122_),
    .ZN(_02123_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05545_ (.I0(\u_cpu.rf_ram.memory[96][6] ),
    .I1(\u_cpu.rf_ram.memory[97][6] ),
    .I2(\u_cpu.rf_ram.memory[98][6] ),
    .I3(\u_cpu.rf_ram.memory[99][6] ),
    .S0(_01567_),
    .S1(_01568_),
    .Z(_02124_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05546_ (.A1(_01548_),
    .A2(_02124_),
    .B(_01579_),
    .ZN(_02125_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05547_ (.I0(\u_cpu.rf_ram.memory[108][6] ),
    .I1(\u_cpu.rf_ram.memory[109][6] ),
    .I2(\u_cpu.rf_ram.memory[110][6] ),
    .I3(\u_cpu.rf_ram.memory[111][6] ),
    .S0(_01529_),
    .S1(_01500_),
    .Z(_02126_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05548_ (.A1(_01512_),
    .A2(_02126_),
    .ZN(_02127_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05549_ (.I0(\u_cpu.rf_ram.memory[104][6] ),
    .I1(\u_cpu.rf_ram.memory[105][6] ),
    .I2(\u_cpu.rf_ram.memory[106][6] ),
    .I3(\u_cpu.rf_ram.memory[107][6] ),
    .S0(_01555_),
    .S1(_01531_),
    .Z(_02128_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05550_ (.A1(_01566_),
    .A2(_02128_),
    .B(_01480_),
    .ZN(_02129_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _05551_ (.A1(_02123_),
    .A2(_02125_),
    .B1(_02127_),
    .B2(_02129_),
    .C(_01560_),
    .ZN(_02130_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05552_ (.I0(\u_cpu.rf_ram.memory[124][6] ),
    .I1(\u_cpu.rf_ram.memory[125][6] ),
    .I2(\u_cpu.rf_ram.memory[126][6] ),
    .I3(\u_cpu.rf_ram.memory[127][6] ),
    .S0(_01496_),
    .S1(_01594_),
    .Z(_02131_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05553_ (.A1(_01543_),
    .A2(_02131_),
    .ZN(_02132_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05554_ (.I0(\u_cpu.rf_ram.memory[120][6] ),
    .I1(\u_cpu.rf_ram.memory[121][6] ),
    .I2(\u_cpu.rf_ram.memory[122][6] ),
    .I3(\u_cpu.rf_ram.memory[123][6] ),
    .S0(_01598_),
    .S1(_01556_),
    .Z(_02133_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05555_ (.A1(_01566_),
    .A2(_02133_),
    .B(_01558_),
    .ZN(_02134_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05556_ (.I0(\u_cpu.rf_ram.memory[112][6] ),
    .I1(\u_cpu.rf_ram.memory[113][6] ),
    .I2(\u_cpu.rf_ram.memory[114][6] ),
    .I3(\u_cpu.rf_ram.memory[115][6] ),
    .S0(_01572_),
    .S1(_01573_),
    .Z(_02135_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05557_ (.A1(_01602_),
    .A2(_02135_),
    .ZN(_02136_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05558_ (.I0(\u_cpu.rf_ram.memory[116][6] ),
    .I1(\u_cpu.rf_ram.memory[117][6] ),
    .I2(\u_cpu.rf_ram.memory[118][6] ),
    .I3(\u_cpu.rf_ram.memory[119][6] ),
    .S0(_01576_),
    .S1(_01577_),
    .Z(_02137_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05559_ (.A1(_01554_),
    .A2(_02137_),
    .B(_01607_),
    .ZN(_02138_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _05560_ (.A1(_02132_),
    .A2(_02134_),
    .B1(_02136_),
    .B2(_02138_),
    .C(_01581_),
    .ZN(_02139_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _05561_ (.A1(_01490_),
    .A2(_02130_),
    .A3(_02139_),
    .ZN(_02140_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05562_ (.I0(\u_cpu.rf_ram.memory[92][6] ),
    .I1(\u_cpu.rf_ram.memory[93][6] ),
    .I2(\u_cpu.rf_ram.memory[94][6] ),
    .I3(\u_cpu.rf_ram.memory[95][6] ),
    .S0(_01562_),
    .S1(_01563_),
    .Z(_02141_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05563_ (.A1(_01464_),
    .A2(_02141_),
    .ZN(_02142_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05564_ (.I0(\u_cpu.rf_ram.memory[88][6] ),
    .I1(\u_cpu.rf_ram.memory[89][6] ),
    .I2(\u_cpu.rf_ram.memory[90][6] ),
    .I3(\u_cpu.rf_ram.memory[91][6] ),
    .S0(_01598_),
    .S1(_01556_),
    .Z(_02143_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05565_ (.A1(_01597_),
    .A2(_02143_),
    .B(_01600_),
    .ZN(_02144_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05566_ (.I0(\u_cpu.rf_ram.memory[80][6] ),
    .I1(\u_cpu.rf_ram.memory[81][6] ),
    .I2(\u_cpu.rf_ram.memory[82][6] ),
    .I3(\u_cpu.rf_ram.memory[83][6] ),
    .S0(_01544_),
    .S1(_01545_),
    .Z(_02145_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05567_ (.A1(_01602_),
    .A2(_02145_),
    .ZN(_02146_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05568_ (.I0(\u_cpu.rf_ram.memory[84][6] ),
    .I1(\u_cpu.rf_ram.memory[85][6] ),
    .I2(\u_cpu.rf_ram.memory[86][6] ),
    .I3(\u_cpu.rf_ram.memory[87][6] ),
    .S0(_01507_),
    .S1(_01605_),
    .Z(_02147_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05569_ (.A1(_01554_),
    .A2(_02147_),
    .B(_01607_),
    .ZN(_02148_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _05570_ (.A1(_02142_),
    .A2(_02144_),
    .B1(_02146_),
    .B2(_02148_),
    .C(_01486_),
    .ZN(_02149_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05571_ (.I0(\u_cpu.rf_ram.memory[64][6] ),
    .I1(\u_cpu.rf_ram.memory[65][6] ),
    .I2(\u_cpu.rf_ram.memory[66][6] ),
    .I3(\u_cpu.rf_ram.memory[67][6] ),
    .S0(_01522_),
    .S1(_01622_),
    .Z(_02150_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05572_ (.A1(_01621_),
    .A2(_02150_),
    .ZN(_02151_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05573_ (.I0(\u_cpu.rf_ram.memory[68][6] ),
    .I1(\u_cpu.rf_ram.memory[69][6] ),
    .I2(\u_cpu.rf_ram.memory[70][6] ),
    .I3(\u_cpu.rf_ram.memory[71][6] ),
    .S0(_01507_),
    .S1(_01605_),
    .Z(_02152_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05574_ (.A1(_01617_),
    .A2(_02152_),
    .B(_01519_),
    .ZN(_02153_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05575_ (.I0(\u_cpu.rf_ram.memory[72][6] ),
    .I1(\u_cpu.rf_ram.memory[73][6] ),
    .I2(\u_cpu.rf_ram.memory[74][6] ),
    .I3(\u_cpu.rf_ram.memory[75][6] ),
    .S0(_01562_),
    .S1(_01563_),
    .Z(_02154_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05576_ (.A1(_01621_),
    .A2(_02154_),
    .ZN(_02155_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05577_ (.I0(\u_cpu.rf_ram.memory[76][6] ),
    .I1(\u_cpu.rf_ram.memory[77][6] ),
    .I2(\u_cpu.rf_ram.memory[78][6] ),
    .I3(\u_cpu.rf_ram.memory[79][6] ),
    .S0(_01529_),
    .S1(_01500_),
    .Z(_02156_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05578_ (.A1(_01617_),
    .A2(_02156_),
    .B(_01600_),
    .ZN(_02157_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _05579_ (.A1(_02151_),
    .A2(_02153_),
    .B1(_02155_),
    .B2(_02157_),
    .C(_01541_),
    .ZN(_02158_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _05580_ (.A1(_01492_),
    .A2(_02149_),
    .A3(_02158_),
    .ZN(_02159_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05581_ (.A1(_02140_),
    .A2(_02159_),
    .B(_01471_),
    .ZN(_02160_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05582_ (.I0(\u_cpu.rf_ram.memory[128][6] ),
    .I1(\u_cpu.rf_ram.memory[129][6] ),
    .I2(\u_cpu.rf_ram.memory[130][6] ),
    .I3(\u_cpu.rf_ram.memory[131][6] ),
    .S0(_01641_),
    .S1(_01635_),
    .Z(_02161_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05583_ (.A1(_01465_),
    .A2(_02161_),
    .ZN(_02162_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05584_ (.I0(\u_cpu.rf_ram.memory[132][6] ),
    .I1(\u_cpu.rf_ram.memory[133][6] ),
    .I2(\u_cpu.rf_ram.memory[134][6] ),
    .I3(\u_cpu.rf_ram.memory[135][6] ),
    .S0(_01634_),
    .S1(_01635_),
    .Z(_02163_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05585_ (.A1(_01638_),
    .A2(_02163_),
    .B(_01482_),
    .ZN(_02164_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05586_ (.I0(\u_cpu.rf_ram.memory[136][6] ),
    .I1(\u_cpu.rf_ram.memory[137][6] ),
    .I2(\u_cpu.rf_ram.memory[138][6] ),
    .I3(\u_cpu.rf_ram.memory[139][6] ),
    .S0(_01523_),
    .S1(_01642_),
    .Z(_02165_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05587_ (.A1(_01493_),
    .A2(_02165_),
    .ZN(_02166_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05588_ (.I0(\u_cpu.rf_ram.memory[140][6] ),
    .I1(\u_cpu.rf_ram.memory[141][6] ),
    .I2(\u_cpu.rf_ram.memory[142][6] ),
    .I3(\u_cpu.rf_ram.memory[143][6] ),
    .S0(_01641_),
    .S1(_01642_),
    .Z(_02167_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05589_ (.A1(_01638_),
    .A2(_02167_),
    .B(_01534_),
    .ZN(_02168_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _05590_ (.A1(_02162_),
    .A2(_02164_),
    .B1(_02166_),
    .B2(_02168_),
    .C(_01466_),
    .ZN(_02169_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05591_ (.A1(_02160_),
    .A2(_02169_),
    .ZN(_02170_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05592_ (.A1(_01473_),
    .A2(_02121_),
    .B(_02170_),
    .ZN(_00006_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05593_ (.I0(\u_cpu.rf_ram.memory[28][7] ),
    .I1(\u_cpu.rf_ram.memory[29][7] ),
    .I2(\u_cpu.rf_ram.memory[30][7] ),
    .I3(\u_cpu.rf_ram.memory[31][7] ),
    .S0(_01497_),
    .S1(_01501_),
    .Z(_02171_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05594_ (.A1(_01513_),
    .A2(_02171_),
    .ZN(_02172_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05595_ (.I0(\u_cpu.rf_ram.memory[24][7] ),
    .I1(\u_cpu.rf_ram.memory[25][7] ),
    .I2(\u_cpu.rf_ram.memory[26][7] ),
    .I3(\u_cpu.rf_ram.memory[27][7] ),
    .S0(_01522_),
    .S1(_01622_),
    .Z(_02173_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05596_ (.A1(_01506_),
    .A2(_02173_),
    .B(_01481_),
    .ZN(_02174_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05597_ (.I0(\u_cpu.rf_ram.memory[20][7] ),
    .I1(\u_cpu.rf_ram.memory[21][7] ),
    .I2(\u_cpu.rf_ram.memory[22][7] ),
    .I3(\u_cpu.rf_ram.memory[23][7] ),
    .S0(_01530_),
    .S1(_01532_),
    .Z(_02175_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05598_ (.A1(_01513_),
    .A2(_02175_),
    .ZN(_02176_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05599_ (.I0(\u_cpu.rf_ram.memory[16][7] ),
    .I1(\u_cpu.rf_ram.memory[17][7] ),
    .I2(\u_cpu.rf_ram.memory[18][7] ),
    .I3(\u_cpu.rf_ram.memory[19][7] ),
    .S0(_01508_),
    .S1(_01509_),
    .Z(_02177_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05600_ (.A1(_01506_),
    .A2(_02177_),
    .B(_01519_),
    .ZN(_02178_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _05601_ (.A1(_02172_),
    .A2(_02174_),
    .B1(_02176_),
    .B2(_02178_),
    .C(_01486_),
    .ZN(_02179_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05602_ (.I0(\u_cpu.rf_ram.memory[4][7] ),
    .I1(\u_cpu.rf_ram.memory[5][7] ),
    .I2(\u_cpu.rf_ram.memory[6][7] ),
    .I3(\u_cpu.rf_ram.memory[7][7] ),
    .S0(_01523_),
    .S1(_01525_),
    .Z(_02180_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05603_ (.A1(_01493_),
    .A2(_02180_),
    .ZN(_02181_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05604_ (.I0(\u_cpu.rf_ram.memory[0][7] ),
    .I1(\u_cpu.rf_ram.memory[1][7] ),
    .I2(\u_cpu.rf_ram.memory[2][7] ),
    .I3(\u_cpu.rf_ram.memory[3][7] ),
    .S0(_01508_),
    .S1(_01509_),
    .Z(_02182_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05605_ (.A1(_01528_),
    .A2(_02182_),
    .B(_01534_),
    .ZN(_02183_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05606_ (.I0(\u_cpu.rf_ram.memory[8][7] ),
    .I1(\u_cpu.rf_ram.memory[9][7] ),
    .I2(\u_cpu.rf_ram.memory[10][7] ),
    .I3(\u_cpu.rf_ram.memory[11][7] ),
    .S0(_01497_),
    .S1(_01501_),
    .Z(_02184_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05607_ (.A1(_01528_),
    .A2(_02184_),
    .ZN(_02185_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05608_ (.I0(\u_cpu.rf_ram.memory[12][7] ),
    .I1(\u_cpu.rf_ram.memory[13][7] ),
    .I2(\u_cpu.rf_ram.memory[14][7] ),
    .I3(\u_cpu.rf_ram.memory[15][7] ),
    .S0(_01530_),
    .S1(_01532_),
    .Z(_02186_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05609_ (.A1(_01464_),
    .A2(_02186_),
    .B(_01481_),
    .ZN(_02187_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _05610_ (.A1(_02181_),
    .A2(_02183_),
    .B1(_02185_),
    .B2(_02187_),
    .C(_01541_),
    .ZN(_02188_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05611_ (.I0(\u_cpu.rf_ram.memory[36][7] ),
    .I1(\u_cpu.rf_ram.memory[37][7] ),
    .I2(\u_cpu.rf_ram.memory[38][7] ),
    .I3(\u_cpu.rf_ram.memory[39][7] ),
    .S0(_01544_),
    .S1(_01545_),
    .Z(_02189_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05612_ (.A1(_01571_),
    .A2(_02189_),
    .ZN(_02190_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05613_ (.I0(\u_cpu.rf_ram.memory[32][7] ),
    .I1(\u_cpu.rf_ram.memory[33][7] ),
    .I2(\u_cpu.rf_ram.memory[34][7] ),
    .I3(\u_cpu.rf_ram.memory[35][7] ),
    .S0(_01495_),
    .S1(_01499_),
    .Z(_02191_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05614_ (.A1(_01504_),
    .A2(_02191_),
    .B(_01518_),
    .ZN(_02192_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05615_ (.I0(\u_cpu.rf_ram.memory[40][7] ),
    .I1(\u_cpu.rf_ram.memory[41][7] ),
    .I2(\u_cpu.rf_ram.memory[42][7] ),
    .I3(\u_cpu.rf_ram.memory[43][7] ),
    .S0(_01551_),
    .S1(_01524_),
    .Z(_02193_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05616_ (.A1(_01505_),
    .A2(_02193_),
    .ZN(_02194_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05617_ (.I0(\u_cpu.rf_ram.memory[44][7] ),
    .I1(\u_cpu.rf_ram.memory[45][7] ),
    .I2(\u_cpu.rf_ram.memory[46][7] ),
    .I3(\u_cpu.rf_ram.memory[47][7] ),
    .S0(_01555_),
    .S1(_01531_),
    .Z(_02195_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05618_ (.A1(_01463_),
    .A2(_02195_),
    .B(_01558_),
    .ZN(_02196_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _05619_ (.A1(_02190_),
    .A2(_02192_),
    .B1(_02194_),
    .B2(_02196_),
    .C(_01560_),
    .ZN(_02197_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05620_ (.I0(\u_cpu.rf_ram.memory[60][7] ),
    .I1(\u_cpu.rf_ram.memory[61][7] ),
    .I2(\u_cpu.rf_ram.memory[62][7] ),
    .I3(\u_cpu.rf_ram.memory[63][7] ),
    .S0(_01496_),
    .S1(_01594_),
    .Z(_02198_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05621_ (.A1(_01543_),
    .A2(_02198_),
    .ZN(_02199_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05622_ (.I0(\u_cpu.rf_ram.memory[56][7] ),
    .I1(\u_cpu.rf_ram.memory[57][7] ),
    .I2(\u_cpu.rf_ram.memory[58][7] ),
    .I3(\u_cpu.rf_ram.memory[59][7] ),
    .S0(_01567_),
    .S1(_01568_),
    .Z(_02200_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05623_ (.A1(_01548_),
    .A2(_02200_),
    .B(_01480_),
    .ZN(_02201_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05624_ (.I0(\u_cpu.rf_ram.memory[52][7] ),
    .I1(\u_cpu.rf_ram.memory[53][7] ),
    .I2(\u_cpu.rf_ram.memory[54][7] ),
    .I3(\u_cpu.rf_ram.memory[55][7] ),
    .S0(_01572_),
    .S1(_01573_),
    .Z(_02202_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05625_ (.A1(_01571_),
    .A2(_02202_),
    .ZN(_02203_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05626_ (.I0(\u_cpu.rf_ram.memory[48][7] ),
    .I1(\u_cpu.rf_ram.memory[49][7] ),
    .I2(\u_cpu.rf_ram.memory[50][7] ),
    .I3(\u_cpu.rf_ram.memory[51][7] ),
    .S0(_01576_),
    .S1(_01577_),
    .Z(_02204_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05627_ (.A1(_01597_),
    .A2(_02204_),
    .B(_01579_),
    .ZN(_02205_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _05628_ (.A1(_02199_),
    .A2(_02201_),
    .B1(_02203_),
    .B2(_02205_),
    .C(_01485_),
    .ZN(_02206_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _05629_ (.A1(_01489_),
    .A2(_02197_),
    .A3(_02206_),
    .Z(_02207_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _05630_ (.A1(_01492_),
    .A2(_02179_),
    .A3(_02188_),
    .B(_02207_),
    .ZN(_02208_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05631_ (.I0(\u_cpu.rf_ram.memory[100][7] ),
    .I1(\u_cpu.rf_ram.memory[101][7] ),
    .I2(\u_cpu.rf_ram.memory[102][7] ),
    .I3(\u_cpu.rf_ram.memory[103][7] ),
    .S0(_01551_),
    .S1(_01524_),
    .Z(_02209_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05632_ (.A1(_01512_),
    .A2(_02209_),
    .ZN(_02210_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05633_ (.I0(\u_cpu.rf_ram.memory[96][7] ),
    .I1(\u_cpu.rf_ram.memory[97][7] ),
    .I2(\u_cpu.rf_ram.memory[98][7] ),
    .I3(\u_cpu.rf_ram.memory[99][7] ),
    .S0(_01567_),
    .S1(_01568_),
    .Z(_02211_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05634_ (.A1(_01548_),
    .A2(_02211_),
    .B(_01518_),
    .ZN(_02212_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05635_ (.I0(\u_cpu.rf_ram.memory[108][7] ),
    .I1(\u_cpu.rf_ram.memory[109][7] ),
    .I2(\u_cpu.rf_ram.memory[110][7] ),
    .I3(\u_cpu.rf_ram.memory[111][7] ),
    .S0(_01529_),
    .S1(_01500_),
    .Z(_02213_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05636_ (.A1(_01512_),
    .A2(_02213_),
    .ZN(_02214_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05637_ (.I0(\u_cpu.rf_ram.memory[104][7] ),
    .I1(\u_cpu.rf_ram.memory[105][7] ),
    .I2(\u_cpu.rf_ram.memory[106][7] ),
    .I3(\u_cpu.rf_ram.memory[107][7] ),
    .S0(_01555_),
    .S1(_01531_),
    .Z(_02215_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05638_ (.A1(_01566_),
    .A2(_02215_),
    .B(_01480_),
    .ZN(_02216_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _05639_ (.A1(_02210_),
    .A2(_02212_),
    .B1(_02214_),
    .B2(_02216_),
    .C(_01560_),
    .ZN(_02217_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05640_ (.I0(\u_cpu.rf_ram.memory[124][7] ),
    .I1(\u_cpu.rf_ram.memory[125][7] ),
    .I2(\u_cpu.rf_ram.memory[126][7] ),
    .I3(\u_cpu.rf_ram.memory[127][7] ),
    .S0(_01496_),
    .S1(_01594_),
    .Z(_02218_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05641_ (.A1(_01543_),
    .A2(_02218_),
    .ZN(_02219_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05642_ (.I0(\u_cpu.rf_ram.memory[120][7] ),
    .I1(\u_cpu.rf_ram.memory[121][7] ),
    .I2(\u_cpu.rf_ram.memory[122][7] ),
    .I3(\u_cpu.rf_ram.memory[123][7] ),
    .S0(_01598_),
    .S1(_01556_),
    .Z(_02220_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05643_ (.A1(_01566_),
    .A2(_02220_),
    .B(_01558_),
    .ZN(_02221_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05644_ (.I0(\u_cpu.rf_ram.memory[112][7] ),
    .I1(\u_cpu.rf_ram.memory[113][7] ),
    .I2(\u_cpu.rf_ram.memory[114][7] ),
    .I3(\u_cpu.rf_ram.memory[115][7] ),
    .S0(_01572_),
    .S1(_01573_),
    .Z(_02222_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05645_ (.A1(_01505_),
    .A2(_02222_),
    .ZN(_02223_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05646_ (.I0(\u_cpu.rf_ram.memory[116][7] ),
    .I1(\u_cpu.rf_ram.memory[117][7] ),
    .I2(\u_cpu.rf_ram.memory[118][7] ),
    .I3(\u_cpu.rf_ram.memory[119][7] ),
    .S0(_01576_),
    .S1(_01577_),
    .Z(_02224_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05647_ (.A1(_01554_),
    .A2(_02224_),
    .B(_01579_),
    .ZN(_02225_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _05648_ (.A1(_02219_),
    .A2(_02221_),
    .B1(_02223_),
    .B2(_02225_),
    .C(_01581_),
    .ZN(_02226_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _05649_ (.A1(_01490_),
    .A2(_02217_),
    .A3(_02226_),
    .ZN(_02227_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05650_ (.I0(\u_cpu.rf_ram.memory[92][7] ),
    .I1(\u_cpu.rf_ram.memory[93][7] ),
    .I2(\u_cpu.rf_ram.memory[94][7] ),
    .I3(\u_cpu.rf_ram.memory[95][7] ),
    .S0(_01562_),
    .S1(_01563_),
    .Z(_02228_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05651_ (.A1(_01464_),
    .A2(_02228_),
    .ZN(_02229_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05652_ (.I0(\u_cpu.rf_ram.memory[88][7] ),
    .I1(\u_cpu.rf_ram.memory[89][7] ),
    .I2(\u_cpu.rf_ram.memory[90][7] ),
    .I3(\u_cpu.rf_ram.memory[91][7] ),
    .S0(_01598_),
    .S1(_01556_),
    .Z(_02230_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05653_ (.A1(_01597_),
    .A2(_02230_),
    .B(_01600_),
    .ZN(_02231_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05654_ (.I0(\u_cpu.rf_ram.memory[80][7] ),
    .I1(\u_cpu.rf_ram.memory[81][7] ),
    .I2(\u_cpu.rf_ram.memory[82][7] ),
    .I3(\u_cpu.rf_ram.memory[83][7] ),
    .S0(_01544_),
    .S1(_01545_),
    .Z(_02232_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05655_ (.A1(_01602_),
    .A2(_02232_),
    .ZN(_02233_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05656_ (.I0(\u_cpu.rf_ram.memory[84][7] ),
    .I1(\u_cpu.rf_ram.memory[85][7] ),
    .I2(\u_cpu.rf_ram.memory[86][7] ),
    .I3(\u_cpu.rf_ram.memory[87][7] ),
    .S0(_01507_),
    .S1(_01605_),
    .Z(_02234_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05657_ (.A1(_01554_),
    .A2(_02234_),
    .B(_01607_),
    .ZN(_02235_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _05658_ (.A1(_02229_),
    .A2(_02231_),
    .B1(_02233_),
    .B2(_02235_),
    .C(_01581_),
    .ZN(_02236_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05659_ (.I0(\u_cpu.rf_ram.memory[64][7] ),
    .I1(\u_cpu.rf_ram.memory[65][7] ),
    .I2(\u_cpu.rf_ram.memory[66][7] ),
    .I3(\u_cpu.rf_ram.memory[67][7] ),
    .S0(_01522_),
    .S1(_01622_),
    .Z(_02237_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05660_ (.A1(_01621_),
    .A2(_02237_),
    .ZN(_02238_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05661_ (.I0(\u_cpu.rf_ram.memory[68][7] ),
    .I1(\u_cpu.rf_ram.memory[69][7] ),
    .I2(\u_cpu.rf_ram.memory[70][7] ),
    .I3(\u_cpu.rf_ram.memory[71][7] ),
    .S0(_01507_),
    .S1(_01605_),
    .Z(_02239_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05662_ (.A1(_01617_),
    .A2(_02239_),
    .B(_01607_),
    .ZN(_02240_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05663_ (.I0(\u_cpu.rf_ram.memory[72][7] ),
    .I1(\u_cpu.rf_ram.memory[73][7] ),
    .I2(\u_cpu.rf_ram.memory[74][7] ),
    .I3(\u_cpu.rf_ram.memory[75][7] ),
    .S0(_01562_),
    .S1(_01563_),
    .Z(_02241_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05664_ (.A1(_01602_),
    .A2(_02241_),
    .ZN(_02242_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05665_ (.I0(\u_cpu.rf_ram.memory[76][7] ),
    .I1(\u_cpu.rf_ram.memory[77][7] ),
    .I2(\u_cpu.rf_ram.memory[78][7] ),
    .I3(\u_cpu.rf_ram.memory[79][7] ),
    .S0(_01529_),
    .S1(_01500_),
    .Z(_02243_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05666_ (.A1(_01617_),
    .A2(_02243_),
    .B(_01600_),
    .ZN(_02244_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _05667_ (.A1(_02238_),
    .A2(_02240_),
    .B1(_02242_),
    .B2(_02244_),
    .C(_01541_),
    .ZN(_02245_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _05668_ (.A1(_01492_),
    .A2(_02236_),
    .A3(_02245_),
    .ZN(_02246_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05669_ (.A1(_02227_),
    .A2(_02246_),
    .B(_01471_),
    .ZN(_02247_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05670_ (.I0(\u_cpu.rf_ram.memory[128][7] ),
    .I1(\u_cpu.rf_ram.memory[129][7] ),
    .I2(\u_cpu.rf_ram.memory[130][7] ),
    .I3(\u_cpu.rf_ram.memory[131][7] ),
    .S0(_01641_),
    .S1(_01642_),
    .Z(_02248_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05671_ (.A1(_01465_),
    .A2(_02248_),
    .ZN(_02249_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05672_ (.I0(\u_cpu.rf_ram.memory[132][7] ),
    .I1(\u_cpu.rf_ram.memory[133][7] ),
    .I2(\u_cpu.rf_ram.memory[134][7] ),
    .I3(\u_cpu.rf_ram.memory[135][7] ),
    .S0(_01634_),
    .S1(_01635_),
    .Z(_02250_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05673_ (.A1(_01638_),
    .A2(_02250_),
    .B(_01482_),
    .ZN(_02251_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05674_ (.I0(\u_cpu.rf_ram.memory[140][7] ),
    .I1(\u_cpu.rf_ram.memory[141][7] ),
    .I2(\u_cpu.rf_ram.memory[142][7] ),
    .I3(\u_cpu.rf_ram.memory[143][7] ),
    .S0(_01523_),
    .S1(_01525_),
    .Z(_02252_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05675_ (.A1(_01638_),
    .A2(_02252_),
    .ZN(_02253_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05676_ (.I0(\u_cpu.rf_ram.memory[136][7] ),
    .I1(\u_cpu.rf_ram.memory[137][7] ),
    .I2(\u_cpu.rf_ram.memory[138][7] ),
    .I3(\u_cpu.rf_ram.memory[139][7] ),
    .S0(_01641_),
    .S1(_01642_),
    .Z(_02254_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05677_ (.A1(_01465_),
    .A2(_02254_),
    .B(_01534_),
    .ZN(_02255_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _05678_ (.A1(_02249_),
    .A2(_02251_),
    .B1(_02253_),
    .B2(_02255_),
    .C(_01466_),
    .ZN(_02256_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05679_ (.A1(_02247_),
    .A2(_02256_),
    .ZN(_02257_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05680_ (.A1(_01473_),
    .A2(_02208_),
    .B(_02257_),
    .ZN(_00007_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _05681_ (.A1(\u_cpu.cpu.state.o_cnt_r[1] ),
    .A2(\u_cpu.cpu.state.o_cnt_r[0] ),
    .A3(\u_cpu.cpu.state.o_cnt_r[3] ),
    .A4(\u_cpu.cpu.state.o_cnt_r[2] ),
    .Z(_02258_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05682_ (.I(_02258_),
    .Z(_02259_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _05683_ (.A1(_01441_),
    .A2(\u_cpu.cpu.bne_or_bge ),
    .Z(_02260_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _05684_ (.A1(\u_arbiter.i_wb_cpu_dbus_we ),
    .A2(\u_cpu.cpu.bufreg.i_sh_signed ),
    .B(_02260_),
    .C(_01445_),
    .ZN(_02261_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05685_ (.A1(\u_cpu.cpu.alu.i_rs1 ),
    .A2(\u_cpu.cpu.alu.add_cy_r ),
    .ZN(_02262_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05686_ (.I(\u_cpu.cpu.bufreg2.i_cnt_done ),
    .Z(_02263_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05687_ (.I(\u_cpu.cpu.immdec.imm11_7[0] ),
    .ZN(_02264_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05688_ (.I(\u_cpu.cpu.decode.opcode[0] ),
    .Z(_02265_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _05689_ (.A1(_01444_),
    .A2(_02265_),
    .A3(\u_cpu.cpu.decode.opcode[1] ),
    .ZN(_02266_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _05690_ (.A1(\u_arbiter.i_wb_cpu_dbus_we ),
    .A2(_02264_),
    .A3(_02266_),
    .Z(_02267_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05691_ (.A1(\u_arbiter.i_wb_cpu_dbus_we ),
    .A2(_02266_),
    .B(\u_cpu.cpu.immdec.imm24_20[0] ),
    .ZN(_02268_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _05692_ (.A1(_01444_),
    .A2(_01445_),
    .A3(_01442_),
    .ZN(_02269_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _05693_ (.A1(_02263_),
    .A2(\u_cpu.cpu.immdec.imm31 ),
    .A3(_02269_),
    .ZN(_02270_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _05694_ (.A1(_02263_),
    .A2(_02267_),
    .A3(_02268_),
    .B(_02270_),
    .ZN(_02271_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05695_ (.I(\u_cpu.rf_ram_if.rtrig1 ),
    .Z(_02272_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _05696_ (.I(\u_cpu.rf_ram.regzero ),
    .ZN(_02273_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05697_ (.A1(\u_cpu.rf_ram.rdata[0] ),
    .A2(_02273_),
    .ZN(_02274_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05698_ (.A1(\u_cpu.rf_ram_if.rdata1[0] ),
    .A2(_02272_),
    .ZN(_02275_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05699_ (.A1(_02272_),
    .A2(_02274_),
    .B(_02275_),
    .ZN(_02276_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05700_ (.I0(_02271_),
    .I1(_02276_),
    .S(\u_arbiter.i_wb_cpu_dbus_we ),
    .Z(_02277_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _05701_ (.A1(_02261_),
    .A2(_02277_),
    .Z(_02278_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05702_ (.A1(\u_cpu.cpu.alu.i_rs1 ),
    .A2(\u_cpu.cpu.alu.add_cy_r ),
    .ZN(_02279_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05703_ (.A1(_02262_),
    .A2(_02278_),
    .B(_02279_),
    .ZN(_02280_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05704_ (.A1(_02259_),
    .A2(_02280_),
    .ZN(_02281_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05705_ (.A1(_02259_),
    .A2(_02261_),
    .B(_02281_),
    .ZN(_00021_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05706_ (.A1(_01441_),
    .A2(\u_cpu.cpu.bne_or_bge ),
    .ZN(_02282_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05707_ (.A1(_01442_),
    .A2(_01439_),
    .ZN(_02283_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05708_ (.A1(_01442_),
    .A2(\u_cpu.cpu.alu.i_rs1 ),
    .B(_02283_),
    .ZN(_02284_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05709_ (.I(_01441_),
    .ZN(_02285_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05710_ (.I(\u_cpu.cpu.bne_or_bge ),
    .ZN(_02286_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05711_ (.A1(_02285_),
    .A2(_02286_),
    .ZN(_02287_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05712_ (.A1(_01441_),
    .A2(_02284_),
    .B(_02286_),
    .ZN(_02288_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05713_ (.A1(_01447_),
    .A2(_01449_),
    .ZN(_02289_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05714_ (.I(\u_cpu.cpu.decode.op22 ),
    .ZN(_02290_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05715_ (.I(\u_cpu.cpu.mem_bytecnt[0] ),
    .Z(_02291_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _05716_ (.A1(\u_cpu.cpu.mem_bytecnt[1] ),
    .A2(\u_cpu.cpu.state.o_cnt[2] ),
    .A3(_02291_),
    .ZN(_02292_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05717_ (.A1(\u_cpu.cpu.decode.op26 ),
    .A2(_01447_),
    .ZN(_02293_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _05718_ (.A1(\u_cpu.cpu.state.o_cnt_r[3] ),
    .A2(_02290_),
    .A3(_02292_),
    .A4(_02293_),
    .Z(_02294_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05719_ (.I(\u_cpu.cpu.genblk3.csr.mcause3_0[0] ),
    .ZN(_02295_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05720_ (.A1(_02263_),
    .A2(\u_cpu.cpu.genblk3.csr.mcause31 ),
    .B(_02292_),
    .ZN(_02296_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _05721_ (.A1(_01448_),
    .A2(\u_cpu.cpu.decode.co_ebreak ),
    .A3(_01447_),
    .ZN(_02297_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05722_ (.A1(_02259_),
    .A2(_02297_),
    .ZN(_02298_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _05723_ (.A1(_02295_),
    .A2(_02292_),
    .B(_02296_),
    .C(_02298_),
    .ZN(_02299_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _05724_ (.A1(_02289_),
    .A2(_02276_),
    .B1(_02294_),
    .B2(\u_cpu.cpu.genblk3.csr.mstatus_mie ),
    .C(_02299_),
    .ZN(_02300_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _05725_ (.A1(_02282_),
    .A2(_02284_),
    .A3(_02287_),
    .B1(_02288_),
    .B2(_02300_),
    .ZN(_02301_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05726_ (.A1(_01460_),
    .A2(_02301_),
    .ZN(_02302_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _05727_ (.A1(\u_cpu.cpu.state.genblk1.misalign_trap_sync_r ),
    .A2(_01459_),
    .Z(_02303_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05728_ (.A1(\u_arbiter.i_wb_cpu_ibus_adr[0] ),
    .A2(_02303_),
    .ZN(_02304_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05729_ (.A1(_02302_),
    .A2(_02304_),
    .ZN(\u_cpu.cpu.o_wdata1 ));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05730_ (.I(_01445_),
    .Z(_02305_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05731_ (.I(\u_cpu.cpu.bufreg.lsb[0] ),
    .Z(_02306_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05732_ (.A1(\u_cpu.cpu.genblk3.csr.o_new_irq ),
    .A2(\u_cpu.cpu.state.init_done ),
    .ZN(_02307_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _05733_ (.A1(_01445_),
    .A2(_02303_),
    .A3(_02307_),
    .ZN(_02308_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05734_ (.I(_01442_),
    .ZN(_02309_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05735_ (.A1(_02285_),
    .A2(_02309_),
    .B(_02260_),
    .ZN(_02310_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _05736_ (.A1(_01445_),
    .A2(_02265_),
    .A3(_02310_),
    .B(_01444_),
    .ZN(_02311_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05737_ (.A1(_02259_),
    .A2(_02311_),
    .ZN(_02312_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05738_ (.I(_01444_),
    .ZN(_02313_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05739_ (.A1(_02313_),
    .A2(_01441_),
    .ZN(_02314_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _05740_ (.A1(_01442_),
    .A2(\u_arbiter.i_wb_cpu_dbus_dat[5] ),
    .B(_02314_),
    .C(\u_cpu.cpu.state.init_done ),
    .ZN(_02315_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _05741_ (.A1(_02308_),
    .A2(_02312_),
    .B1(_02315_),
    .B2(\u_cpu.cpu.state.stage_two_req ),
    .ZN(_02316_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _05742_ (.A1(_02306_),
    .A2(_02316_),
    .Z(_02317_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05743_ (.A1(_01444_),
    .A2(_02265_),
    .ZN(_02318_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05744_ (.A1(_01445_),
    .A2(_02318_),
    .ZN(_02319_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _05745_ (.A1(\u_cpu.cpu.immdec.imm31 ),
    .A2(_02269_),
    .Z(_02320_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _05746_ (.A1(_02263_),
    .A2(_02267_),
    .A3(_02268_),
    .ZN(_02321_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05747_ (.A1(_02263_),
    .A2(_02320_),
    .B(_02321_),
    .ZN(_02322_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05748_ (.A1(\u_cpu.cpu.state.o_cnt[2] ),
    .A2(_02291_),
    .B(\u_cpu.cpu.mem_bytecnt[1] ),
    .ZN(_02323_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05749_ (.A1(_02322_),
    .A2(_02323_),
    .B(_02319_),
    .ZN(_02324_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05750_ (.I(\u_cpu.cpu.decode.co_ebreak ),
    .ZN(_02325_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _05751_ (.A1(_01445_),
    .A2(\u_arbiter.i_wb_cpu_dbus_we ),
    .B1(_02325_),
    .B2(_01457_),
    .ZN(_02326_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05752_ (.I(_02265_),
    .ZN(_02327_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05753_ (.I(\u_cpu.cpu.decode.opcode[1] ),
    .ZN(_02328_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05754_ (.A1(_02327_),
    .A2(_02328_),
    .ZN(_02329_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _05755_ (.A1(_02266_),
    .A2(_02326_),
    .A3(_02329_),
    .B(\u_arbiter.i_wb_cpu_ibus_adr[0] ),
    .ZN(_02330_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05756_ (.I(_02330_),
    .ZN(_02331_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _05757_ (.A1(\u_cpu.cpu.ctrl.pc_plus_offset_cy_r ),
    .A2(_02331_),
    .Z(_02332_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _05758_ (.A1(_02317_),
    .A2(_02319_),
    .B(_02324_),
    .C(_02332_),
    .ZN(_02333_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05759_ (.A1(\u_cpu.cpu.state.o_cnt_r[0] ),
    .A2(_02292_),
    .ZN(_02334_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05760_ (.I(_02316_),
    .Z(_02335_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05761_ (.A1(_02306_),
    .A2(_02335_),
    .ZN(_02336_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05762_ (.A1(_02322_),
    .A2(_02323_),
    .ZN(_02337_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05763_ (.A1(_02319_),
    .A2(_02337_),
    .ZN(_02338_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _05764_ (.A1(\u_cpu.cpu.ctrl.pc_plus_offset_cy_r ),
    .A2(_02330_),
    .Z(_02339_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _05765_ (.A1(_02336_),
    .A2(_02319_),
    .B(_02338_),
    .C(_02339_),
    .ZN(_02340_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _05766_ (.A1(_02333_),
    .A2(_02334_),
    .A3(_02340_),
    .ZN(_02341_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05767_ (.A1(_02305_),
    .A2(_02317_),
    .ZN(_02342_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05768_ (.A1(_02305_),
    .A2(_02341_),
    .B(_02342_),
    .ZN(_02343_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05769_ (.A1(\u_cpu.cpu.alu.i_rs1 ),
    .A2(_02277_),
    .ZN(_02344_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05770_ (.A1(_01441_),
    .A2(_02344_),
    .ZN(_02345_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05771_ (.A1(\u_cpu.cpu.alu.i_rs1 ),
    .A2(_02277_),
    .B(_01442_),
    .ZN(_02346_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _05772_ (.A1(\u_cpu.cpu.bne_or_bge ),
    .A2(_02344_),
    .B(_02345_),
    .C(_02346_),
    .ZN(_02347_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _05773_ (.A1(\u_cpu.cpu.alu.i_rs1 ),
    .A2(\u_cpu.cpu.alu.add_cy_r ),
    .A3(_02278_),
    .Z(_02348_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _05774_ (.A1(_01441_),
    .A2(_02309_),
    .A3(\u_cpu.cpu.alu.cmp_r ),
    .ZN(_02349_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _05775_ (.A1(_01443_),
    .A2(_02348_),
    .B1(_02349_),
    .B2(_02334_),
    .C(_02336_),
    .ZN(_02350_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05776_ (.A1(_02347_),
    .A2(_02350_),
    .ZN(_02351_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _05777_ (.A1(_02313_),
    .A2(_02305_),
    .A3(_02265_),
    .A4(_02351_),
    .ZN(_02352_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05778_ (.I(\u_cpu.cpu.mem_if.signbit ),
    .ZN(_02353_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _05779_ (.A1(_02285_),
    .A2(\u_cpu.cpu.mem_bytecnt[1] ),
    .B1(_02291_),
    .B2(_02282_),
    .ZN(_02354_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05780_ (.I(\u_cpu.cpu.bufreg.lsb[1] ),
    .Z(_02355_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05781_ (.I0(\u_arbiter.i_wb_cpu_dbus_dat[0] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_dat[8] ),
    .I2(\u_arbiter.i_wb_cpu_dbus_dat[16] ),
    .I3(\u_arbiter.i_wb_cpu_dbus_dat[24] ),
    .S0(_02306_),
    .S1(_02355_),
    .Z(_02356_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05782_ (.A1(_02354_),
    .A2(_02356_),
    .ZN(_02357_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05783_ (.A1(_02353_),
    .A2(_02354_),
    .B(_02357_),
    .ZN(_00798_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _05784_ (.A1(_01442_),
    .A2(_02357_),
    .B(_01444_),
    .C(_02265_),
    .ZN(_02358_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05785_ (.I(\u_cpu.cpu.state.o_cnt_r[1] ),
    .ZN(_02359_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05786_ (.A1(_02359_),
    .A2(\u_cpu.cpu.ctrl.i_iscomp ),
    .ZN(_02360_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _05787_ (.A1(\u_cpu.cpu.state.o_cnt_r[2] ),
    .A2(\u_cpu.cpu.ctrl.i_iscomp ),
    .B(_02292_),
    .C(_02360_),
    .ZN(_02361_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _05788_ (.A1(\u_cpu.cpu.ctrl.pc_plus_4_cy_r ),
    .A2(\u_arbiter.i_wb_cpu_ibus_adr[0] ),
    .Z(_02362_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _05789_ (.A1(_02361_),
    .A2(_02362_),
    .Z(_02363_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05790_ (.A1(_01445_),
    .A2(_02265_),
    .ZN(_02364_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _05791_ (.A1(_02363_),
    .A2(_02364_),
    .B(_01460_),
    .C(_02300_),
    .ZN(_02365_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05792_ (.A1(_00798_),
    .A2(_02358_),
    .B(_02365_),
    .ZN(_02366_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _05793_ (.A1(_02305_),
    .A2(_02318_),
    .A3(_02341_),
    .B(_02366_),
    .ZN(_02367_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _05794_ (.A1(_01460_),
    .A2(_02343_),
    .B1(_02352_),
    .B2(_02367_),
    .ZN(_02368_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _05795_ (.I(_02368_),
    .ZN(\u_cpu.cpu.o_wdata0 ));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05796_ (.A1(_02273_),
    .A2(\u_cpu.rf_ram.rdata[1] ),
    .ZN(_02369_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05797_ (.A1(_02272_),
    .A2(\u_cpu.rf_ram_if.rdata1[1] ),
    .ZN(_02370_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05798_ (.A1(_02272_),
    .A2(_02369_),
    .B(_02370_),
    .ZN(_00015_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05799_ (.A1(_02273_),
    .A2(\u_cpu.rf_ram.rdata[2] ),
    .ZN(_02371_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05800_ (.A1(_02272_),
    .A2(\u_cpu.rf_ram_if.rdata1[2] ),
    .ZN(_02372_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05801_ (.A1(_02272_),
    .A2(_02371_),
    .B(_02372_),
    .ZN(_00016_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05802_ (.A1(_02273_),
    .A2(\u_cpu.rf_ram.rdata[3] ),
    .ZN(_02373_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05803_ (.A1(_02272_),
    .A2(\u_cpu.rf_ram_if.rdata1[3] ),
    .ZN(_02374_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05804_ (.A1(_02272_),
    .A2(_02373_),
    .B(_02374_),
    .ZN(_00017_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05805_ (.A1(_02273_),
    .A2(\u_cpu.rf_ram.rdata[4] ),
    .ZN(_02375_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05806_ (.A1(_02272_),
    .A2(\u_cpu.rf_ram_if.rdata1[4] ),
    .ZN(_02376_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05807_ (.A1(_02272_),
    .A2(_02375_),
    .B(_02376_),
    .ZN(_00018_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05808_ (.A1(_02273_),
    .A2(\u_cpu.rf_ram.rdata[5] ),
    .ZN(_02377_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05809_ (.A1(_02272_),
    .A2(\u_cpu.rf_ram_if.rdata1[5] ),
    .ZN(_02378_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05810_ (.A1(_02272_),
    .A2(_02377_),
    .B(_02378_),
    .ZN(_00019_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05811_ (.A1(_02273_),
    .A2(\u_cpu.rf_ram.rdata[6] ),
    .ZN(_02379_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05812_ (.A1(_02272_),
    .A2(\u_cpu.rf_ram_if.rdata1[6] ),
    .ZN(_02380_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05813_ (.A1(_02272_),
    .A2(_02379_),
    .B(_02380_),
    .ZN(_00020_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05814_ (.A1(\u_cpu.rf_ram_if.rdata0[1] ),
    .A2(_01467_),
    .ZN(_02381_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05815_ (.A1(_01467_),
    .A2(_02274_),
    .B(_02381_),
    .ZN(_00008_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05816_ (.A1(\u_cpu.rf_ram_if.rdata0[2] ),
    .A2(_01467_),
    .ZN(_02382_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05817_ (.A1(_01467_),
    .A2(_02369_),
    .B(_02382_),
    .ZN(_00009_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05818_ (.A1(\u_cpu.rf_ram_if.rdata0[3] ),
    .A2(_01467_),
    .ZN(_02383_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05819_ (.A1(_01467_),
    .A2(_02371_),
    .B(_02383_),
    .ZN(_00010_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05820_ (.A1(\u_cpu.rf_ram_if.rdata0[4] ),
    .A2(_01467_),
    .ZN(_02384_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05821_ (.A1(_01467_),
    .A2(_02373_),
    .B(_02384_),
    .ZN(_00011_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05822_ (.A1(\u_cpu.rf_ram_if.rdata0[5] ),
    .A2(_01467_),
    .ZN(_02385_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05823_ (.A1(_01467_),
    .A2(_02375_),
    .B(_02385_),
    .ZN(_00012_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05824_ (.A1(\u_cpu.rf_ram_if.rdata0[6] ),
    .A2(_01467_),
    .ZN(_02386_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05825_ (.A1(_01467_),
    .A2(_02377_),
    .B(_02386_),
    .ZN(_00013_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05826_ (.A1(\u_cpu.rf_ram_if.rdata0[7] ),
    .A2(_01467_),
    .ZN(_02387_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05827_ (.A1(_01467_),
    .A2(_02379_),
    .B(_02387_),
    .ZN(_00014_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05828_ (.I(io_in[3]),
    .Z(_02388_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05829_ (.I(_02388_),
    .Z(_02389_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05830_ (.A1(io_in[2]),
    .A2(_02389_),
    .ZN(_02390_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _05831_ (.A1(_01441_),
    .A2(_02355_),
    .B1(_02260_),
    .B2(_02306_),
    .ZN(_02391_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _05832_ (.A1(\u_cpu.cpu.state.o_cnt_r[1] ),
    .A2(\u_cpu.cpu.state.o_cnt_r[0] ),
    .A3(\u_cpu.cpu.state.o_cnt_r[3] ),
    .A4(\u_cpu.cpu.state.o_cnt_r[2] ),
    .ZN(_02392_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05833_ (.A1(\u_cpu.cpu.state.init_done ),
    .A2(_02392_),
    .ZN(_02393_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _05834_ (.A1(_01444_),
    .A2(_02305_),
    .A3(_02393_),
    .ZN(_02394_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05835_ (.I(io_in[1]),
    .Z(_02395_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05836_ (.I(_02395_),
    .ZN(_02396_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05837_ (.A1(_02396_),
    .A2(\u_cpu.cpu.state.ibus_cyc ),
    .ZN(_02397_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05838_ (.A1(_02388_),
    .A2(_02397_),
    .ZN(_02398_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05839_ (.A1(_02391_),
    .A2(_02394_),
    .B(_02398_),
    .ZN(_02399_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05840_ (.A1(_02390_),
    .A2(_02399_),
    .ZN(_00026_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05841_ (.I(\u_arbiter.i_wb_cpu_dbus_we ),
    .ZN(_02400_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05842_ (.I(_02388_),
    .ZN(_02401_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05843_ (.I(_02401_),
    .Z(_02402_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05844_ (.I(_02402_),
    .Z(_02403_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05845_ (.A1(_02403_),
    .A2(\u_cpu.cpu.genblk3.csr.i_mtip ),
    .ZN(_02404_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05846_ (.A1(_02400_),
    .A2(_02398_),
    .B(_02404_),
    .ZN(_00037_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05847_ (.A1(_02306_),
    .A2(_02355_),
    .B(_02388_),
    .ZN(_02405_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05848_ (.A1(\u_arbiter.i_wb_cpu_ack ),
    .A2(_02389_),
    .B(_02405_),
    .ZN(_02406_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _05849_ (.I(_02406_),
    .ZN(_00048_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05850_ (.A1(\u_cpu.cpu.bne_or_bge ),
    .A2(_02306_),
    .ZN(_02407_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05851_ (.A1(_01441_),
    .A2(_02402_),
    .ZN(_02408_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05852_ (.A1(_02355_),
    .A2(_02407_),
    .B(_02408_),
    .ZN(_02409_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05853_ (.A1(\u_arbiter.i_wb_cpu_rdt[0] ),
    .A2(_02389_),
    .B(_02409_),
    .ZN(_02410_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _05854_ (.I(_02410_),
    .ZN(_00059_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05855_ (.I(\u_arbiter.i_wb_cpu_rdt[1] ),
    .ZN(_02411_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05856_ (.I(_02306_),
    .ZN(_02412_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05857_ (.A1(_02412_),
    .A2(_02355_),
    .ZN(_02413_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _05858_ (.A1(_02411_),
    .A2(_02403_),
    .B1(_02413_),
    .B2(_02408_),
    .ZN(_00070_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05859_ (.I(\u_arbiter.i_wb_cpu_rdt[2] ),
    .ZN(_02414_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05860_ (.A1(\u_cpu.cpu.bne_or_bge ),
    .A2(_02306_),
    .B(_02355_),
    .ZN(_02415_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _05861_ (.A1(_02414_),
    .A2(_02403_),
    .B1(_02408_),
    .B2(_02415_),
    .ZN(_00081_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05862_ (.I(\u_arbiter.i_wb_cpu_rdt[3] ),
    .ZN(_02416_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05863_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[0] ),
    .A2(_02389_),
    .ZN(_02417_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05864_ (.A1(_02416_),
    .A2(_02389_),
    .B(_02417_),
    .ZN(_00092_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05865_ (.I(_02388_),
    .Z(_02418_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05866_ (.I0(\u_arbiter.i_wb_cpu_rdt[4] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_dat[1] ),
    .S(_02418_),
    .Z(_02419_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05867_ (.I(_02419_),
    .Z(_00093_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05868_ (.I0(\u_arbiter.i_wb_cpu_rdt[5] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_dat[2] ),
    .S(_02418_),
    .Z(_02420_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05869_ (.I(_02420_),
    .Z(_00094_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05870_ (.I0(\u_arbiter.i_wb_cpu_rdt[6] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_dat[3] ),
    .S(_02418_),
    .Z(_02421_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05871_ (.I(_02421_),
    .Z(_00095_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05872_ (.I0(\u_arbiter.i_wb_cpu_rdt[7] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_dat[4] ),
    .S(_02418_),
    .Z(_02422_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05873_ (.I(_02422_),
    .Z(_00027_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05874_ (.I0(\u_arbiter.i_wb_cpu_rdt[8] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_dat[5] ),
    .S(_02418_),
    .Z(_02423_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05875_ (.I(_02423_),
    .Z(_00028_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05876_ (.I0(\u_arbiter.i_wb_cpu_rdt[9] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_dat[6] ),
    .S(_02418_),
    .Z(_02424_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05877_ (.I(_02424_),
    .Z(_00029_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05878_ (.I0(\u_arbiter.i_wb_cpu_rdt[10] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_dat[7] ),
    .S(_02418_),
    .Z(_02425_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05879_ (.I(_02425_),
    .Z(_00030_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05880_ (.I0(\u_arbiter.i_wb_cpu_rdt[11] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_dat[8] ),
    .S(_02418_),
    .Z(_02426_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05881_ (.I(_02426_),
    .Z(_00031_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05882_ (.I0(\u_arbiter.i_wb_cpu_rdt[12] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_dat[9] ),
    .S(_02418_),
    .Z(_02427_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05883_ (.I(_02427_),
    .Z(_00032_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05884_ (.I0(\u_arbiter.i_wb_cpu_rdt[13] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_dat[10] ),
    .S(_02418_),
    .Z(_02428_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05885_ (.I(_02428_),
    .Z(_00033_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05886_ (.I0(\u_arbiter.i_wb_cpu_rdt[14] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_dat[11] ),
    .S(_02418_),
    .Z(_02429_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05887_ (.I(_02429_),
    .Z(_00034_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05888_ (.I0(\u_arbiter.i_wb_cpu_rdt[15] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_dat[12] ),
    .S(_02418_),
    .Z(_02430_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05889_ (.I(_02430_),
    .Z(_00035_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05890_ (.I(_02388_),
    .Z(_02431_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05891_ (.I0(\u_arbiter.i_wb_cpu_rdt[16] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_dat[13] ),
    .S(_02431_),
    .Z(_02432_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05892_ (.I(_02432_),
    .Z(_00036_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05893_ (.I0(\u_arbiter.i_wb_cpu_rdt[17] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_dat[14] ),
    .S(_02431_),
    .Z(_02433_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05894_ (.I(_02433_),
    .Z(_00038_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05895_ (.I0(\u_arbiter.i_wb_cpu_rdt[18] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_dat[15] ),
    .S(_02431_),
    .Z(_02434_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05896_ (.I(_02434_),
    .Z(_00039_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05897_ (.I0(\u_arbiter.i_wb_cpu_rdt[19] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_dat[16] ),
    .S(_02431_),
    .Z(_02435_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05898_ (.I(_02435_),
    .Z(_00040_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05899_ (.I0(\u_arbiter.i_wb_cpu_rdt[20] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_dat[17] ),
    .S(_02431_),
    .Z(_02436_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05900_ (.I(_02436_),
    .Z(_00041_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05901_ (.I0(\u_arbiter.i_wb_cpu_rdt[21] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_dat[18] ),
    .S(_02431_),
    .Z(_02437_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05902_ (.I(_02437_),
    .Z(_00042_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05903_ (.I0(\u_arbiter.i_wb_cpu_rdt[22] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_dat[19] ),
    .S(_02431_),
    .Z(_02438_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05904_ (.I(_02438_),
    .Z(_00043_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05905_ (.I0(\u_arbiter.i_wb_cpu_rdt[23] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_dat[20] ),
    .S(_02431_),
    .Z(_02439_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05906_ (.I(_02439_),
    .Z(_00044_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05907_ (.I0(\u_arbiter.i_wb_cpu_rdt[24] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_dat[21] ),
    .S(_02431_),
    .Z(_02440_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05908_ (.I(_02440_),
    .Z(_00045_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05909_ (.I0(\u_arbiter.i_wb_cpu_rdt[25] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_dat[22] ),
    .S(_02431_),
    .Z(_02441_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05910_ (.I(_02441_),
    .Z(_00046_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05911_ (.I0(\u_arbiter.i_wb_cpu_rdt[26] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_dat[23] ),
    .S(_02431_),
    .Z(_02442_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05912_ (.I(_02442_),
    .Z(_00047_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05913_ (.I0(\u_arbiter.i_wb_cpu_rdt[27] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_dat[24] ),
    .S(_02431_),
    .Z(_02443_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05914_ (.I(_02443_),
    .Z(_00049_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05915_ (.I0(\u_arbiter.i_wb_cpu_rdt[28] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_dat[25] ),
    .S(_02431_),
    .Z(_02444_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05916_ (.I(_02444_),
    .Z(_00050_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05917_ (.I(\u_arbiter.i_wb_cpu_dbus_dat[26] ),
    .ZN(_02445_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05918_ (.A1(\u_arbiter.i_wb_cpu_rdt[29] ),
    .A2(_02403_),
    .ZN(_02446_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05919_ (.A1(_02445_),
    .A2(_02403_),
    .B(_02446_),
    .ZN(_00051_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05920_ (.I0(\u_arbiter.i_wb_cpu_rdt[30] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_dat[27] ),
    .S(_02431_),
    .Z(_02447_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05921_ (.I(_02447_),
    .Z(_00052_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05922_ (.I0(\u_arbiter.i_wb_cpu_rdt[31] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_dat[28] ),
    .S(_02431_),
    .Z(_02448_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05923_ (.I(_02448_),
    .Z(_00053_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05924_ (.I0(\u_scanchain_local.module_data_in[34] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_dat[29] ),
    .S(_02431_),
    .Z(_02449_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05925_ (.I(_02449_),
    .Z(_00054_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05926_ (.I(\u_arbiter.i_wb_cpu_dbus_dat[30] ),
    .ZN(_02450_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05927_ (.A1(_02403_),
    .A2(\u_scanchain_local.module_data_in[35] ),
    .ZN(_02451_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05928_ (.A1(_02450_),
    .A2(_02403_),
    .B(_02451_),
    .ZN(_00055_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05929_ (.I(\u_arbiter.i_wb_cpu_dbus_dat[31] ),
    .ZN(_02452_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05930_ (.A1(_02403_),
    .A2(\u_scanchain_local.module_data_in[36] ),
    .ZN(_02453_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05931_ (.A1(_02452_),
    .A2(_02403_),
    .B(_02453_),
    .ZN(_00056_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05932_ (.A1(_02403_),
    .A2(\u_scanchain_local.module_data_in[37] ),
    .ZN(_02454_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05933_ (.A1(_02401_),
    .A2(_02397_),
    .ZN(_02455_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05934_ (.I(_02455_),
    .Z(_02456_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05935_ (.A1(\u_arbiter.i_wb_cpu_ibus_adr[0] ),
    .A2(_02456_),
    .ZN(_02457_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05936_ (.A1(_02454_),
    .A2(_02457_),
    .ZN(_00057_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05937_ (.A1(_02403_),
    .A2(\u_scanchain_local.module_data_in[38] ),
    .ZN(_02458_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05938_ (.A1(\u_arbiter.i_wb_cpu_ibus_adr[1] ),
    .A2(_02456_),
    .ZN(_02459_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05939_ (.A1(_02458_),
    .A2(_02459_),
    .ZN(_00058_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _05940_ (.A1(_02396_),
    .A2(\u_cpu.cpu.state.ibus_cyc ),
    .Z(_02460_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05941_ (.I(_02460_),
    .Z(_02461_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05942_ (.A1(_02388_),
    .A2(_02461_),
    .ZN(_02462_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05943_ (.I(_02462_),
    .Z(_02463_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05944_ (.I(\u_cpu.cpu.genblk1.align.ctrl_misal ),
    .Z(_02464_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05945_ (.I(_02464_),
    .Z(_02465_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05946_ (.I(_02465_),
    .Z(_02466_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05947_ (.I(_02466_),
    .Z(_02467_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _05948_ (.A1(_02467_),
    .A2(\u_cpu.cpu.ctrl.o_ibus_adr[2] ),
    .Z(_02468_));
 gf180mcu_fd_sc_mcu7t5v0__oai222_1 _05949_ (.A1(_02389_),
    .A2(\u_scanchain_local.module_data_in[39] ),
    .B1(_02463_),
    .B2(_02468_),
    .C1(_02398_),
    .C2(\u_arbiter.i_wb_cpu_dbus_adr[2] ),
    .ZN(_02469_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _05950_ (.I(_02469_),
    .ZN(_00060_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05951_ (.A1(_02467_),
    .A2(\u_cpu.cpu.ctrl.o_ibus_adr[2] ),
    .ZN(_02470_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _05952_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[3] ),
    .A2(_02470_),
    .Z(_02471_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _05953_ (.A1(_02389_),
    .A2(\u_scanchain_local.module_data_in[40] ),
    .B1(_02398_),
    .B2(\u_arbiter.i_wb_cpu_dbus_adr[3] ),
    .ZN(_02472_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05954_ (.A1(_02456_),
    .A2(_02471_),
    .B(_02472_),
    .ZN(_00061_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _05955_ (.A1(_02467_),
    .A2(\u_cpu.cpu.ctrl.o_ibus_adr[3] ),
    .A3(\u_cpu.cpu.ctrl.o_ibus_adr[2] ),
    .ZN(_02473_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _05956_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[4] ),
    .A2(_02473_),
    .Z(_02474_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _05957_ (.A1(_02389_),
    .A2(\u_scanchain_local.module_data_in[41] ),
    .B1(_02398_),
    .B2(\u_arbiter.i_wb_cpu_dbus_adr[4] ),
    .ZN(_02475_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05958_ (.A1(_02456_),
    .A2(_02474_),
    .B(_02475_),
    .ZN(_00062_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _05959_ (.A1(_02464_),
    .A2(\u_cpu.cpu.ctrl.o_ibus_adr[4] ),
    .A3(\u_cpu.cpu.ctrl.o_ibus_adr[3] ),
    .A4(\u_cpu.cpu.ctrl.o_ibus_adr[2] ),
    .Z(_02476_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _05960_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[5] ),
    .A2(_02476_),
    .ZN(_02477_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05961_ (.A1(_02401_),
    .A2(_02461_),
    .ZN(_02478_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _05962_ (.A1(_02403_),
    .A2(\u_scanchain_local.module_data_in[42] ),
    .B1(_02478_),
    .B2(\u_arbiter.i_wb_cpu_dbus_adr[5] ),
    .ZN(_02479_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05963_ (.A1(_02463_),
    .A2(_02477_),
    .B(_02479_),
    .ZN(_00063_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05964_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[5] ),
    .A2(_02476_),
    .ZN(_02480_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _05965_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[6] ),
    .A2(_02480_),
    .Z(_02481_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _05966_ (.A1(_02418_),
    .A2(\u_scanchain_local.module_data_in[43] ),
    .B1(_02398_),
    .B2(\u_arbiter.i_wb_cpu_dbus_adr[6] ),
    .ZN(_02482_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05967_ (.A1(_02456_),
    .A2(_02481_),
    .B(_02482_),
    .ZN(_00064_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _05968_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[6] ),
    .A2(\u_cpu.cpu.ctrl.o_ibus_adr[5] ),
    .A3(_02476_),
    .ZN(_02483_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _05969_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[7] ),
    .A2(_02483_),
    .Z(_02484_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _05970_ (.A1(_02418_),
    .A2(\u_scanchain_local.module_data_in[44] ),
    .B1(_02398_),
    .B2(\u_arbiter.i_wb_cpu_dbus_adr[7] ),
    .ZN(_02485_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05971_ (.A1(_02456_),
    .A2(_02484_),
    .B(_02485_),
    .ZN(_00065_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05972_ (.I(\u_cpu.cpu.ctrl.o_ibus_adr[8] ),
    .ZN(_02486_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _05973_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[7] ),
    .A2(\u_cpu.cpu.ctrl.o_ibus_adr[6] ),
    .A3(\u_cpu.cpu.ctrl.o_ibus_adr[5] ),
    .A4(_02476_),
    .ZN(_02487_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05974_ (.A1(_02486_),
    .A2(_02487_),
    .ZN(_02488_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05975_ (.A1(_02486_),
    .A2(_02487_),
    .ZN(_02489_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05976_ (.A1(_02456_),
    .A2(_02489_),
    .ZN(_02490_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _05977_ (.A1(_02403_),
    .A2(\u_scanchain_local.module_data_in[45] ),
    .B1(_02478_),
    .B2(\u_arbiter.i_wb_cpu_dbus_adr[8] ),
    .ZN(_02491_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05978_ (.A1(_02488_),
    .A2(_02490_),
    .B(_02491_),
    .ZN(_00066_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05979_ (.I(\u_cpu.cpu.ctrl.o_ibus_adr[9] ),
    .ZN(_02492_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _05980_ (.A1(_02492_),
    .A2(_02486_),
    .A3(_02487_),
    .ZN(_02493_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05981_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[9] ),
    .A2(_02488_),
    .B(_02456_),
    .ZN(_02494_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _05982_ (.A1(_02403_),
    .A2(\u_scanchain_local.module_data_in[46] ),
    .B1(_02478_),
    .B2(\u_arbiter.i_wb_cpu_dbus_adr[9] ),
    .ZN(_02495_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05983_ (.A1(_02493_),
    .A2(_02494_),
    .B(_02495_),
    .ZN(_00067_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _05984_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[10] ),
    .A2(_02493_),
    .ZN(_02496_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _05985_ (.A1(_02403_),
    .A2(\u_scanchain_local.module_data_in[47] ),
    .B1(_02478_),
    .B2(\u_arbiter.i_wb_cpu_dbus_adr[10] ),
    .ZN(_02497_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05986_ (.A1(_02463_),
    .A2(_02496_),
    .B(_02497_),
    .ZN(_00068_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05987_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[11] ),
    .A2(\u_cpu.cpu.ctrl.o_ibus_adr[10] ),
    .ZN(_02498_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _05988_ (.A1(_02492_),
    .A2(_02486_),
    .A3(_02487_),
    .A4(_02498_),
    .ZN(_02499_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05989_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[10] ),
    .A2(_02493_),
    .B(\u_cpu.cpu.ctrl.o_ibus_adr[11] ),
    .ZN(_02500_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05990_ (.A1(_02499_),
    .A2(_02500_),
    .B(_02456_),
    .ZN(_02501_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _05991_ (.A1(_02389_),
    .A2(\u_scanchain_local.module_data_in[48] ),
    .B1(_02398_),
    .B2(\u_arbiter.i_wb_cpu_dbus_adr[11] ),
    .C(_02501_),
    .ZN(_02502_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _05992_ (.I(_02502_),
    .ZN(_00069_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05993_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[12] ),
    .A2(_02499_),
    .B(_02461_),
    .ZN(_02503_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05994_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[12] ),
    .A2(_02499_),
    .B(_02503_),
    .ZN(_02504_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05995_ (.A1(\u_arbiter.i_wb_cpu_dbus_adr[12] ),
    .A2(_02397_),
    .B(_02504_),
    .ZN(_02505_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05996_ (.A1(_02389_),
    .A2(\u_scanchain_local.module_data_in[49] ),
    .ZN(_02506_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05997_ (.A1(_02389_),
    .A2(_02505_),
    .B(_02506_),
    .ZN(_00071_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05998_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[12] ),
    .A2(_02499_),
    .B(\u_cpu.cpu.ctrl.o_ibus_adr[13] ),
    .ZN(_02507_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _05999_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[13] ),
    .A2(\u_cpu.cpu.ctrl.o_ibus_adr[12] ),
    .A3(_02499_),
    .Z(_02508_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06000_ (.A1(_02402_),
    .A2(\u_scanchain_local.module_data_in[50] ),
    .B1(_02478_),
    .B2(\u_arbiter.i_wb_cpu_dbus_adr[13] ),
    .ZN(_02509_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _06001_ (.A1(_02463_),
    .A2(_02507_),
    .A3(_02508_),
    .B(_02509_),
    .ZN(_00072_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _06002_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[14] ),
    .A2(_02508_),
    .ZN(_02510_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06003_ (.A1(_02402_),
    .A2(\u_scanchain_local.module_data_in[51] ),
    .B1(_02478_),
    .B2(\u_arbiter.i_wb_cpu_dbus_adr[14] ),
    .ZN(_02511_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06004_ (.A1(_02463_),
    .A2(_02510_),
    .B(_02511_),
    .ZN(_00073_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06005_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[14] ),
    .A2(_02508_),
    .ZN(_02512_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06006_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[15] ),
    .A2(_02512_),
    .Z(_02513_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _06007_ (.A1(_02418_),
    .A2(\u_scanchain_local.module_data_in[52] ),
    .B1(_02398_),
    .B2(\u_arbiter.i_wb_cpu_dbus_adr[15] ),
    .ZN(_02514_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06008_ (.A1(_02456_),
    .A2(_02513_),
    .B(_02514_),
    .ZN(_00074_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06009_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[15] ),
    .A2(\u_cpu.cpu.ctrl.o_ibus_adr[14] ),
    .A3(_02508_),
    .ZN(_02515_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06010_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[16] ),
    .A2(_02515_),
    .Z(_02516_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _06011_ (.A1(_02418_),
    .A2(\u_scanchain_local.module_data_in[53] ),
    .B1(_02398_),
    .B2(\u_arbiter.i_wb_cpu_dbus_adr[16] ),
    .ZN(_02517_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06012_ (.A1(_02456_),
    .A2(_02516_),
    .B(_02517_),
    .ZN(_00075_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06013_ (.I(\u_cpu.cpu.ctrl.o_ibus_adr[16] ),
    .ZN(_02518_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06014_ (.A1(_02518_),
    .A2(_02515_),
    .ZN(_02519_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _06015_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[17] ),
    .A2(\u_cpu.cpu.ctrl.o_ibus_adr[16] ),
    .A3(\u_cpu.cpu.ctrl.o_ibus_adr[15] ),
    .A4(\u_cpu.cpu.ctrl.o_ibus_adr[14] ),
    .Z(_02520_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _06016_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[13] ),
    .A2(\u_cpu.cpu.ctrl.o_ibus_adr[12] ),
    .A3(_02499_),
    .A4(_02520_),
    .ZN(_02521_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _06017_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[17] ),
    .A2(_02519_),
    .B(_02521_),
    .C(_02461_),
    .ZN(_02522_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06018_ (.A1(\u_arbiter.i_wb_cpu_dbus_adr[17] ),
    .A2(_02397_),
    .ZN(_02523_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06019_ (.A1(_02388_),
    .A2(_02522_),
    .A3(_02523_),
    .ZN(_02524_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06020_ (.A1(_02389_),
    .A2(\u_scanchain_local.module_data_in[54] ),
    .B(_02524_),
    .ZN(_02525_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _06021_ (.I(_02525_),
    .ZN(_00076_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06022_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[18] ),
    .A2(_02521_),
    .Z(_02526_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06023_ (.A1(_02402_),
    .A2(\u_scanchain_local.module_data_in[55] ),
    .B1(_02478_),
    .B2(\u_arbiter.i_wb_cpu_dbus_adr[18] ),
    .ZN(_02527_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06024_ (.A1(_02463_),
    .A2(_02526_),
    .B(_02527_),
    .ZN(_00077_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06025_ (.I(\u_cpu.cpu.ctrl.o_ibus_adr[18] ),
    .ZN(_02528_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06026_ (.I(\u_cpu.cpu.ctrl.o_ibus_adr[19] ),
    .ZN(_02529_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06027_ (.A1(_02528_),
    .A2(_02521_),
    .B(_02529_),
    .ZN(_02530_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _06028_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[19] ),
    .A2(\u_cpu.cpu.ctrl.o_ibus_adr[18] ),
    .A3(_02508_),
    .A4(_02520_),
    .ZN(_02531_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06029_ (.A1(_02461_),
    .A2(_02530_),
    .A3(_02531_),
    .ZN(_02532_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06030_ (.A1(\u_arbiter.i_wb_cpu_dbus_adr[19] ),
    .A2(_02397_),
    .ZN(_02533_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06031_ (.A1(_02388_),
    .A2(_02532_),
    .A3(_02533_),
    .ZN(_02534_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06032_ (.A1(_02389_),
    .A2(\u_scanchain_local.module_data_in[56] ),
    .B(_02534_),
    .ZN(_02535_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _06033_ (.I(_02535_),
    .ZN(_00078_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06034_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[20] ),
    .A2(_02531_),
    .Z(_02536_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06035_ (.A1(_02402_),
    .A2(\u_scanchain_local.module_data_in[57] ),
    .B1(_02478_),
    .B2(\u_arbiter.i_wb_cpu_dbus_adr[20] ),
    .ZN(_02537_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06036_ (.A1(_02463_),
    .A2(_02536_),
    .B(_02537_),
    .ZN(_00079_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06037_ (.I(\u_cpu.cpu.ctrl.o_ibus_adr[20] ),
    .ZN(_02538_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _06038_ (.A1(_02538_),
    .A2(_02529_),
    .A3(_02528_),
    .A4(_02521_),
    .ZN(_02539_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06039_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[21] ),
    .A2(_02539_),
    .ZN(_02540_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06040_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[21] ),
    .A2(_02539_),
    .ZN(_02541_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06041_ (.A1(_02456_),
    .A2(_02541_),
    .ZN(_02542_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06042_ (.A1(_02402_),
    .A2(\u_scanchain_local.module_data_in[58] ),
    .B1(_02478_),
    .B2(\u_arbiter.i_wb_cpu_dbus_adr[21] ),
    .ZN(_02543_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06043_ (.A1(_02540_),
    .A2(_02542_),
    .B(_02543_),
    .ZN(_00080_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06044_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[22] ),
    .A2(_02541_),
    .Z(_02544_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06045_ (.A1(_02402_),
    .A2(\u_scanchain_local.module_data_in[59] ),
    .B1(_02478_),
    .B2(\u_arbiter.i_wb_cpu_dbus_adr[22] ),
    .ZN(_02545_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06046_ (.A1(_02463_),
    .A2(_02544_),
    .B(_02545_),
    .ZN(_00082_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _06047_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[22] ),
    .A2(\u_cpu.cpu.ctrl.o_ibus_adr[21] ),
    .A3(_02539_),
    .Z(_02546_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06048_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[23] ),
    .A2(_02546_),
    .ZN(_02547_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _06049_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[23] ),
    .A2(\u_cpu.cpu.ctrl.o_ibus_adr[22] ),
    .A3(\u_cpu.cpu.ctrl.o_ibus_adr[21] ),
    .A4(_02539_),
    .ZN(_02548_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06050_ (.A1(_02461_),
    .A2(_02548_),
    .ZN(_02549_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06051_ (.A1(\u_arbiter.i_wb_cpu_dbus_adr[23] ),
    .A2(_02397_),
    .ZN(_02550_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _06052_ (.A1(_02547_),
    .A2(_02549_),
    .B(_02550_),
    .C(_02388_),
    .ZN(_02551_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06053_ (.A1(_02389_),
    .A2(\u_scanchain_local.module_data_in[60] ),
    .B(_02551_),
    .ZN(_02552_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _06054_ (.I(_02552_),
    .ZN(_00083_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06055_ (.A1(_02389_),
    .A2(\u_scanchain_local.module_data_in[61] ),
    .ZN(_02553_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06056_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[24] ),
    .A2(\u_cpu.cpu.ctrl.o_ibus_adr[23] ),
    .A3(_02546_),
    .ZN(_02554_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06057_ (.I(\u_cpu.cpu.ctrl.o_ibus_adr[24] ),
    .ZN(_02555_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06058_ (.A1(_02555_),
    .A2(_02548_),
    .B(_02397_),
    .ZN(_02556_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _06059_ (.A1(\u_arbiter.i_wb_cpu_dbus_adr[24] ),
    .A2(_02397_),
    .B1(_02554_),
    .B2(_02556_),
    .C(_02402_),
    .ZN(_02557_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06060_ (.A1(_02553_),
    .A2(_02557_),
    .ZN(_00084_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06061_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[25] ),
    .A2(_02554_),
    .Z(_02558_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06062_ (.A1(_02402_),
    .A2(\u_scanchain_local.module_data_in[62] ),
    .B1(_02478_),
    .B2(\u_arbiter.i_wb_cpu_dbus_adr[25] ),
    .ZN(_02559_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06063_ (.A1(_02463_),
    .A2(_02558_),
    .B(_02559_),
    .ZN(_00085_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06064_ (.I(\u_cpu.cpu.ctrl.o_ibus_adr[26] ),
    .ZN(_02560_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06065_ (.I(\u_cpu.cpu.ctrl.o_ibus_adr[25] ),
    .ZN(_02561_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _06066_ (.A1(_02560_),
    .A2(_02561_),
    .A3(_02555_),
    .A4(_02548_),
    .ZN(_02562_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06067_ (.A1(_02561_),
    .A2(_02554_),
    .ZN(_02563_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06068_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[26] ),
    .A2(_02563_),
    .B(_02456_),
    .ZN(_02564_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06069_ (.A1(_02402_),
    .A2(\u_scanchain_local.module_data_in[63] ),
    .B1(_02478_),
    .B2(\u_arbiter.i_wb_cpu_dbus_adr[26] ),
    .ZN(_02565_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06070_ (.A1(_02562_),
    .A2(_02564_),
    .B(_02565_),
    .ZN(_00086_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06071_ (.I(\u_scanchain_local.module_data_in[64] ),
    .ZN(_02566_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06072_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[27] ),
    .A2(_02562_),
    .B(_02397_),
    .ZN(_02567_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06073_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[27] ),
    .A2(_02562_),
    .B(_02567_),
    .ZN(_02568_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06074_ (.A1(\u_arbiter.i_wb_cpu_dbus_adr[27] ),
    .A2(_02397_),
    .B(_02402_),
    .ZN(_02569_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06075_ (.A1(_02403_),
    .A2(_02566_),
    .B1(_02568_),
    .B2(_02569_),
    .ZN(_00087_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06076_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[27] ),
    .A2(_02562_),
    .B(\u_cpu.cpu.ctrl.o_ibus_adr[28] ),
    .ZN(_02570_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06077_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[28] ),
    .A2(\u_cpu.cpu.ctrl.o_ibus_adr[27] ),
    .A3(_02562_),
    .ZN(_02571_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06078_ (.A1(_02456_),
    .A2(_02571_),
    .ZN(_02572_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06079_ (.A1(_02402_),
    .A2(\u_scanchain_local.module_data_in[65] ),
    .B1(_02478_),
    .B2(\u_arbiter.i_wb_cpu_dbus_adr[28] ),
    .ZN(_02573_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06080_ (.A1(_02570_),
    .A2(_02572_),
    .B(_02573_),
    .ZN(_00088_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06081_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[29] ),
    .A2(_02571_),
    .Z(_02574_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06082_ (.A1(_02402_),
    .A2(\u_scanchain_local.module_data_in[66] ),
    .B1(_02478_),
    .B2(\u_arbiter.i_wb_cpu_dbus_adr[29] ),
    .ZN(_02575_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06083_ (.A1(_02463_),
    .A2(_02574_),
    .B(_02575_),
    .ZN(_00089_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06084_ (.A1(_02389_),
    .A2(\u_scanchain_local.module_data_in[67] ),
    .ZN(_02576_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _06085_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[29] ),
    .A2(\u_cpu.cpu.ctrl.o_ibus_adr[28] ),
    .A3(\u_cpu.cpu.ctrl.o_ibus_adr[27] ),
    .A4(_02562_),
    .Z(_02577_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06086_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[30] ),
    .A2(_02577_),
    .ZN(_02578_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06087_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[30] ),
    .A2(_02577_),
    .ZN(_02579_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06088_ (.A1(_02397_),
    .A2(_02579_),
    .ZN(_02580_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _06089_ (.A1(\u_arbiter.i_wb_cpu_dbus_adr[30] ),
    .A2(_02397_),
    .B1(_02578_),
    .B2(_02580_),
    .C(_02402_),
    .ZN(_02581_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06090_ (.A1(_02576_),
    .A2(_02581_),
    .ZN(_00090_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06091_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[31] ),
    .A2(_02578_),
    .Z(_02582_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06092_ (.A1(_02402_),
    .A2(\u_scanchain_local.module_data_in[68] ),
    .B1(_02478_),
    .B2(\u_arbiter.i_wb_cpu_dbus_adr[31] ),
    .ZN(_02583_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06093_ (.A1(_02463_),
    .A2(_02582_),
    .B(_02583_),
    .ZN(_00091_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06094_ (.A1(_02305_),
    .A2(\u_cpu.cpu.decode.opcode[1] ),
    .ZN(_02584_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06095_ (.A1(_01445_),
    .A2(_02327_),
    .ZN(_02585_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _06096_ (.A1(\u_cpu.cpu.alu.i_rs1 ),
    .A2(\u_cpu.cpu.bufreg.c_r ),
    .A3(_02584_),
    .A4(_02585_),
    .ZN(_02586_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06097_ (.A1(_02265_),
    .A2(\u_cpu.cpu.decode.opcode[1] ),
    .ZN(_02587_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06098_ (.A1(_02587_),
    .A2(_02329_),
    .B(_02305_),
    .ZN(_02588_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06099_ (.A1(_02334_),
    .A2(_02588_),
    .B(_02313_),
    .ZN(_02589_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06100_ (.A1(_02322_),
    .A2(_02589_),
    .ZN(_02590_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06101_ (.A1(\u_cpu.cpu.alu.i_rs1 ),
    .A2(_02584_),
    .A3(_02585_),
    .ZN(_02591_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _06102_ (.A1(\u_cpu.cpu.bufreg.c_r ),
    .A2(_02591_),
    .ZN(_02592_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06103_ (.A1(_02590_),
    .A2(_02592_),
    .ZN(_02593_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06104_ (.A1(_02308_),
    .A2(_02312_),
    .ZN(_02594_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06105_ (.A1(\u_cpu.cpu.state.stage_two_req ),
    .A2(_02315_),
    .ZN(_02595_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06106_ (.A1(_02594_),
    .A2(_02595_),
    .ZN(_02596_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06107_ (.A1(_02586_),
    .A2(_02593_),
    .B(_02596_),
    .ZN(_00022_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06108_ (.A1(\u_cpu.cpu.ctrl.pc_plus_offset_cy_r ),
    .A2(_02331_),
    .ZN(_02597_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06109_ (.A1(_02307_),
    .A2(_02311_),
    .ZN(_02598_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06110_ (.A1(_02259_),
    .A2(_02598_),
    .ZN(_02599_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06111_ (.A1(_02597_),
    .A2(_02333_),
    .B(_02599_),
    .ZN(_00024_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06112_ (.A1(\u_cpu.cpu.ctrl.pc_plus_4_cy_r ),
    .A2(\u_arbiter.i_wb_cpu_ibus_adr[0] ),
    .ZN(_02600_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06113_ (.I(_02361_),
    .ZN(_02601_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06114_ (.A1(_02601_),
    .A2(_02362_),
    .ZN(_02602_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06115_ (.A1(_02600_),
    .A2(_02602_),
    .B(_02599_),
    .ZN(_00023_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06116_ (.A1(_01460_),
    .A2(_01456_),
    .B(_02392_),
    .ZN(\u_cpu.cpu.o_wen1 ));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _06117_ (.A1(\u_cpu.cpu.immdec.imm11_7[1] ),
    .A2(\u_cpu.cpu.immdec.imm11_7[2] ),
    .A3(\u_cpu.cpu.immdec.imm11_7[3] ),
    .A4(\u_cpu.cpu.immdec.imm11_7[0] ),
    .Z(_02603_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _06118_ (.A1(_02265_),
    .A2(\u_arbiter.i_wb_cpu_dbus_we ),
    .B(_02364_),
    .C(_02313_),
    .ZN(_02604_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _06119_ (.A1(\u_cpu.cpu.immdec.imm11_7[4] ),
    .A2(_02603_),
    .B(_02604_),
    .C(_02598_),
    .ZN(_02605_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06120_ (.A1(_01460_),
    .A2(_02605_),
    .B(_02392_),
    .ZN(\u_cpu.cpu.o_wen0 ));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06121_ (.I(\u_cpu.rf_ram_if.genblk1.wtrig0_r ),
    .Z(_02606_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _06122_ (.A1(_02303_),
    .A2(_01455_),
    .Z(_02607_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06123_ (.A1(_02606_),
    .A2(_02303_),
    .ZN(_02608_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06124_ (.A1(_02606_),
    .A2(_02607_),
    .B1(_02608_),
    .B2(_02264_),
    .ZN(_02609_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06125_ (.A1(\u_cpu.cpu.decode.op26 ),
    .A2(\u_cpu.cpu.decode.co_ebreak ),
    .A3(_02606_),
    .ZN(_02610_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _06126_ (.I(_02606_),
    .ZN(_02611_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06127_ (.A1(\u_cpu.cpu.immdec.imm11_7[1] ),
    .A2(_02611_),
    .ZN(_02612_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06128_ (.A1(_01460_),
    .A2(_02610_),
    .A3(_02612_),
    .ZN(_02613_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _06129_ (.A1(_02609_),
    .A2(_02613_),
    .Z(_02614_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06130_ (.A1(\u_cpu.rf_ram_if.rcnt[0] ),
    .A2(\u_cpu.rf_ram_if.rcnt[1] ),
    .B(\u_cpu.rf_ram_if.rcnt[2] ),
    .ZN(_02615_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06131_ (.A1(_01494_),
    .A2(_02615_),
    .Z(_02616_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06132_ (.I(_02616_),
    .ZN(_02617_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06133_ (.A1(_01500_),
    .A2(_02617_),
    .ZN(_02618_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06134_ (.A1(_02614_),
    .A2(_02618_),
    .ZN(_02619_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06135_ (.A1(\u_cpu.cpu.immdec.imm11_7[2] ),
    .A2(_02608_),
    .ZN(_02620_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06136_ (.I(\u_cpu.cpu.immdec.imm11_7[4] ),
    .ZN(_02621_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06137_ (.A1(_02606_),
    .A2(\u_cpu.rf_ram_if.wen1_r ),
    .B1(\u_cpu.rf_ram_if.rtrig0 ),
    .B2(\u_cpu.rf_ram_if.wen0_r ),
    .ZN(_02622_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06138_ (.A1(_02621_),
    .A2(_02622_),
    .ZN(_02623_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06139_ (.A1(_02608_),
    .A2(_02623_),
    .ZN(_02624_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _06140_ (.A1(\u_cpu.cpu.immdec.imm11_7[3] ),
    .A2(_02620_),
    .A3(_02624_),
    .ZN(_02625_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06141_ (.I(_02625_),
    .Z(_02626_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06142_ (.A1(_02619_),
    .A2(_02626_),
    .ZN(_02627_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06143_ (.I(_02627_),
    .Z(_02628_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06144_ (.A1(\u_cpu.rf_ram_if.wdata1_r[0] ),
    .A2(_02606_),
    .Z(_02629_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06145_ (.A1(\u_cpu.rf_ram_if.wdata0_r[0] ),
    .A2(_02611_),
    .B(_02629_),
    .ZN(_02630_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06146_ (.I(_02630_),
    .Z(_02631_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06147_ (.I(_02631_),
    .Z(_02632_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06148_ (.A1(\u_cpu.rf_ram.memory[82][0] ),
    .A2(_02628_),
    .ZN(_02633_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06149_ (.A1(_02628_),
    .A2(_02632_),
    .B(_02633_),
    .ZN(_00096_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06150_ (.A1(_02606_),
    .A2(\u_cpu.rf_ram_if.wdata1_r[1] ),
    .Z(_02634_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06151_ (.A1(_02611_),
    .A2(\u_cpu.rf_ram_if.wdata0_r[1] ),
    .B(_02634_),
    .ZN(_02635_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06152_ (.I(_02635_),
    .Z(_02636_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06153_ (.I(_02636_),
    .Z(_02637_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06154_ (.A1(\u_cpu.rf_ram.memory[82][1] ),
    .A2(_02628_),
    .ZN(_02638_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06155_ (.A1(_02628_),
    .A2(_02637_),
    .B(_02638_),
    .ZN(_00097_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06156_ (.A1(_02606_),
    .A2(\u_cpu.rf_ram_if.wdata1_r[2] ),
    .Z(_02639_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06157_ (.A1(_02611_),
    .A2(\u_cpu.rf_ram_if.wdata0_r[2] ),
    .B(_02639_),
    .ZN(_02640_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06158_ (.I(_02640_),
    .Z(_02641_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06159_ (.I(_02641_),
    .Z(_02642_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06160_ (.A1(\u_cpu.rf_ram.memory[82][2] ),
    .A2(_02628_),
    .ZN(_02643_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06161_ (.A1(_02628_),
    .A2(_02642_),
    .B(_02643_),
    .ZN(_00098_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06162_ (.A1(_02606_),
    .A2(\u_cpu.rf_ram_if.wdata1_r[3] ),
    .Z(_02644_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06163_ (.A1(_02611_),
    .A2(\u_cpu.rf_ram_if.wdata0_r[3] ),
    .B(_02644_),
    .ZN(_02645_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06164_ (.I(_02645_),
    .Z(_02646_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06165_ (.I(_02646_),
    .Z(_02647_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06166_ (.A1(\u_cpu.rf_ram.memory[82][3] ),
    .A2(_02628_),
    .ZN(_02648_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06167_ (.A1(_02628_),
    .A2(_02647_),
    .B(_02648_),
    .ZN(_00099_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06168_ (.A1(_02606_),
    .A2(\u_cpu.rf_ram_if.wdata1_r[4] ),
    .Z(_02649_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06169_ (.A1(_02611_),
    .A2(\u_cpu.rf_ram_if.wdata0_r[4] ),
    .B(_02649_),
    .ZN(_02650_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06170_ (.I(_02650_),
    .Z(_02651_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06171_ (.I(_02651_),
    .Z(_02652_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06172_ (.A1(\u_cpu.rf_ram.memory[82][4] ),
    .A2(_02628_),
    .ZN(_02653_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06173_ (.A1(_02628_),
    .A2(_02652_),
    .B(_02653_),
    .ZN(_00100_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06174_ (.A1(_02606_),
    .A2(\u_cpu.rf_ram_if.wdata1_r[5] ),
    .Z(_02654_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06175_ (.A1(_02611_),
    .A2(\u_cpu.rf_ram_if.wdata0_r[5] ),
    .B(_02654_),
    .ZN(_02655_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06176_ (.I(_02655_),
    .Z(_02656_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06177_ (.I(_02656_),
    .Z(_02657_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06178_ (.A1(\u_cpu.rf_ram.memory[82][5] ),
    .A2(_02628_),
    .ZN(_02658_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06179_ (.A1(_02628_),
    .A2(_02657_),
    .B(_02658_),
    .ZN(_00101_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06180_ (.A1(_02606_),
    .A2(\u_cpu.rf_ram_if.wdata1_r[6] ),
    .Z(_02659_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06181_ (.A1(_02611_),
    .A2(\u_cpu.rf_ram_if.wdata0_r[6] ),
    .B(_02659_),
    .ZN(_02660_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06182_ (.I(_02660_),
    .Z(_02661_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06183_ (.I(_02661_),
    .Z(_02662_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06184_ (.A1(\u_cpu.rf_ram.memory[82][6] ),
    .A2(_02628_),
    .ZN(_02663_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06185_ (.A1(_02628_),
    .A2(_02662_),
    .B(_02663_),
    .ZN(_00102_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06186_ (.I(\u_cpu.rf_ram_if.wdata1_r[7] ),
    .ZN(_02664_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06187_ (.I0(_02664_),
    .I1(_02368_),
    .S(_02611_),
    .Z(_02665_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06188_ (.I(_02665_),
    .Z(_02666_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06189_ (.I(_02666_),
    .Z(_02667_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06190_ (.A1(\u_cpu.rf_ram.memory[82][7] ),
    .A2(_02628_),
    .ZN(_02668_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06191_ (.A1(_02628_),
    .A2(_02667_),
    .B(_02668_),
    .ZN(_00103_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06192_ (.I(_02631_),
    .Z(_02669_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _06193_ (.A1(\u_cpu.rf_ram_if.rcnt[0] ),
    .A2(\u_cpu.rf_ram_if.rcnt[1] ),
    .B(_01494_),
    .C(\u_cpu.rf_ram_if.rcnt[2] ),
    .ZN(_02670_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06194_ (.A1(_01498_),
    .A2(_02670_),
    .Z(_02671_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _06195_ (.A1(_02617_),
    .A2(_02671_),
    .Z(_02672_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _06196_ (.A1(_01460_),
    .A2(_02610_),
    .A3(_02612_),
    .Z(_02673_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06197_ (.A1(_02609_),
    .A2(_02673_),
    .ZN(_02674_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06198_ (.A1(_02672_),
    .A2(_02674_),
    .ZN(_02675_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _06199_ (.A1(\u_cpu.cpu.immdec.imm11_7[3] ),
    .A2(\u_cpu.cpu.immdec.imm11_7[4] ),
    .A3(_02620_),
    .A4(_02622_),
    .ZN(_02676_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06200_ (.I(_02676_),
    .Z(_02677_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06201_ (.A1(_02675_),
    .A2(_02677_),
    .ZN(_02678_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06202_ (.I(_02678_),
    .Z(_02679_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06203_ (.A1(\u_cpu.rf_ram.memory[21][0] ),
    .A2(_02679_),
    .ZN(_02680_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06204_ (.A1(_02669_),
    .A2(_02679_),
    .B(_02680_),
    .ZN(_00104_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06205_ (.I(_02636_),
    .Z(_02681_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06206_ (.A1(\u_cpu.rf_ram.memory[21][1] ),
    .A2(_02679_),
    .ZN(_02682_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06207_ (.A1(_02681_),
    .A2(_02679_),
    .B(_02682_),
    .ZN(_00105_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06208_ (.I(_02641_),
    .Z(_02683_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06209_ (.A1(\u_cpu.rf_ram.memory[21][2] ),
    .A2(_02679_),
    .ZN(_02684_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06210_ (.A1(_02683_),
    .A2(_02679_),
    .B(_02684_),
    .ZN(_00106_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06211_ (.I(_02646_),
    .Z(_02685_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06212_ (.A1(\u_cpu.rf_ram.memory[21][3] ),
    .A2(_02679_),
    .ZN(_02686_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06213_ (.A1(_02685_),
    .A2(_02679_),
    .B(_02686_),
    .ZN(_00107_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06214_ (.I(_02651_),
    .Z(_02687_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06215_ (.A1(\u_cpu.rf_ram.memory[21][4] ),
    .A2(_02679_),
    .ZN(_02688_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06216_ (.A1(_02687_),
    .A2(_02679_),
    .B(_02688_),
    .ZN(_00108_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06217_ (.I(_02656_),
    .Z(_02689_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06218_ (.A1(\u_cpu.rf_ram.memory[21][5] ),
    .A2(_02679_),
    .ZN(_02690_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06219_ (.A1(_02689_),
    .A2(_02679_),
    .B(_02690_),
    .ZN(_00109_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06220_ (.I(_02661_),
    .Z(_02691_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06221_ (.A1(\u_cpu.rf_ram.memory[21][6] ),
    .A2(_02679_),
    .ZN(_02692_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06222_ (.A1(_02691_),
    .A2(_02679_),
    .B(_02692_),
    .ZN(_00110_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06223_ (.I(_02666_),
    .Z(_02693_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06224_ (.A1(\u_cpu.rf_ram.memory[21][7] ),
    .A2(_02679_),
    .ZN(_02694_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06225_ (.A1(_02693_),
    .A2(_02679_),
    .B(_02694_),
    .ZN(_00111_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06226_ (.A1(_02614_),
    .A2(_02672_),
    .ZN(_02695_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06227_ (.A1(_02626_),
    .A2(_02695_),
    .ZN(_02696_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06228_ (.I(_02696_),
    .Z(_02697_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06229_ (.A1(\u_cpu.rf_ram.memory[81][0] ),
    .A2(_02697_),
    .ZN(_02698_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06230_ (.A1(_02669_),
    .A2(_02697_),
    .B(_02698_),
    .ZN(_00112_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06231_ (.A1(\u_cpu.rf_ram.memory[81][1] ),
    .A2(_02697_),
    .ZN(_02699_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06232_ (.A1(_02681_),
    .A2(_02697_),
    .B(_02699_),
    .ZN(_00113_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06233_ (.A1(\u_cpu.rf_ram.memory[81][2] ),
    .A2(_02697_),
    .ZN(_02700_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06234_ (.A1(_02683_),
    .A2(_02697_),
    .B(_02700_),
    .ZN(_00114_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06235_ (.A1(\u_cpu.rf_ram.memory[81][3] ),
    .A2(_02697_),
    .ZN(_02701_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06236_ (.A1(_02685_),
    .A2(_02697_),
    .B(_02701_),
    .ZN(_00115_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06237_ (.A1(\u_cpu.rf_ram.memory[81][4] ),
    .A2(_02697_),
    .ZN(_02702_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06238_ (.A1(_02687_),
    .A2(_02697_),
    .B(_02702_),
    .ZN(_00116_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06239_ (.A1(\u_cpu.rf_ram.memory[81][5] ),
    .A2(_02697_),
    .ZN(_02703_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06240_ (.A1(_02689_),
    .A2(_02697_),
    .B(_02703_),
    .ZN(_00117_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06241_ (.A1(\u_cpu.rf_ram.memory[81][6] ),
    .A2(_02697_),
    .ZN(_02704_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06242_ (.A1(_02691_),
    .A2(_02697_),
    .B(_02704_),
    .ZN(_00118_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06243_ (.A1(\u_cpu.rf_ram.memory[81][7] ),
    .A2(_02697_),
    .ZN(_02705_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06244_ (.A1(_02693_),
    .A2(_02697_),
    .B(_02705_),
    .ZN(_00119_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06245_ (.A1(_02619_),
    .A2(_02677_),
    .ZN(_02706_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06246_ (.I(_02706_),
    .Z(_02707_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06247_ (.A1(\u_cpu.rf_ram.memory[18][0] ),
    .A2(_02707_),
    .ZN(_02708_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06248_ (.A1(_02669_),
    .A2(_02707_),
    .B(_02708_),
    .ZN(_00120_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06249_ (.A1(\u_cpu.rf_ram.memory[18][1] ),
    .A2(_02707_),
    .ZN(_02709_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06250_ (.A1(_02681_),
    .A2(_02707_),
    .B(_02709_),
    .ZN(_00121_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06251_ (.A1(\u_cpu.rf_ram.memory[18][2] ),
    .A2(_02707_),
    .ZN(_02710_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06252_ (.A1(_02683_),
    .A2(_02707_),
    .B(_02710_),
    .ZN(_00122_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06253_ (.A1(\u_cpu.rf_ram.memory[18][3] ),
    .A2(_02707_),
    .ZN(_02711_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06254_ (.A1(_02685_),
    .A2(_02707_),
    .B(_02711_),
    .ZN(_00123_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06255_ (.A1(\u_cpu.rf_ram.memory[18][4] ),
    .A2(_02707_),
    .ZN(_02712_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06256_ (.A1(_02687_),
    .A2(_02707_),
    .B(_02712_),
    .ZN(_00124_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06257_ (.A1(\u_cpu.rf_ram.memory[18][5] ),
    .A2(_02707_),
    .ZN(_02713_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06258_ (.A1(_02689_),
    .A2(_02707_),
    .B(_02713_),
    .ZN(_00125_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06259_ (.A1(\u_cpu.rf_ram.memory[18][6] ),
    .A2(_02707_),
    .ZN(_02714_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06260_ (.A1(_02691_),
    .A2(_02707_),
    .B(_02714_),
    .ZN(_00126_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06261_ (.A1(\u_cpu.rf_ram.memory[18][7] ),
    .A2(_02707_),
    .ZN(_02715_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06262_ (.A1(_02693_),
    .A2(_02707_),
    .B(_02715_),
    .ZN(_00127_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _06263_ (.A1(_01563_),
    .A2(_02616_),
    .Z(_02716_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06264_ (.A1(_02674_),
    .A2(_02716_),
    .ZN(_02717_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06265_ (.A1(_02677_),
    .A2(_02717_),
    .ZN(_02718_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06266_ (.I(_02718_),
    .Z(_02719_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06267_ (.A1(\u_cpu.rf_ram.memory[20][0] ),
    .A2(_02719_),
    .ZN(_02720_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06268_ (.A1(_02669_),
    .A2(_02719_),
    .B(_02720_),
    .ZN(_00128_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06269_ (.A1(\u_cpu.rf_ram.memory[20][1] ),
    .A2(_02719_),
    .ZN(_02721_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06270_ (.A1(_02681_),
    .A2(_02719_),
    .B(_02721_),
    .ZN(_00129_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06271_ (.A1(\u_cpu.rf_ram.memory[20][2] ),
    .A2(_02719_),
    .ZN(_02722_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06272_ (.A1(_02683_),
    .A2(_02719_),
    .B(_02722_),
    .ZN(_00130_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06273_ (.A1(\u_cpu.rf_ram.memory[20][3] ),
    .A2(_02719_),
    .ZN(_02723_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06274_ (.A1(_02685_),
    .A2(_02719_),
    .B(_02723_),
    .ZN(_00131_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06275_ (.A1(\u_cpu.rf_ram.memory[20][4] ),
    .A2(_02719_),
    .ZN(_02724_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06276_ (.A1(_02687_),
    .A2(_02719_),
    .B(_02724_),
    .ZN(_00132_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06277_ (.A1(\u_cpu.rf_ram.memory[20][5] ),
    .A2(_02719_),
    .ZN(_02725_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06278_ (.A1(_02689_),
    .A2(_02719_),
    .B(_02725_),
    .ZN(_00133_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06279_ (.A1(\u_cpu.rf_ram.memory[20][6] ),
    .A2(_02719_),
    .ZN(_02726_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06280_ (.A1(_02691_),
    .A2(_02719_),
    .B(_02726_),
    .ZN(_00134_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06281_ (.A1(\u_cpu.rf_ram.memory[20][7] ),
    .A2(_02719_),
    .ZN(_02727_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06282_ (.A1(_02693_),
    .A2(_02719_),
    .B(_02727_),
    .ZN(_00135_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06283_ (.I(\u_cpu.cpu.immdec.imm11_7[2] ),
    .ZN(_02728_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06284_ (.A1(\u_cpu.cpu.immdec.imm11_7[3] ),
    .A2(_02608_),
    .ZN(_02729_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06285_ (.A1(_02728_),
    .A2(_02608_),
    .A3(_02729_),
    .ZN(_02730_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _06286_ (.A1(\u_cpu.cpu.immdec.imm11_7[4] ),
    .A2(_02622_),
    .A3(_02730_),
    .ZN(_02731_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06287_ (.A1(_02695_),
    .A2(_02731_),
    .Z(_02732_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06288_ (.I(_02732_),
    .Z(_02733_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06289_ (.A1(\u_cpu.rf_ram.memory[1][0] ),
    .A2(_02733_),
    .ZN(_02734_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06290_ (.A1(_02632_),
    .A2(_02733_),
    .B(_02734_),
    .ZN(_00136_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06291_ (.A1(\u_cpu.rf_ram.memory[1][1] ),
    .A2(_02733_),
    .ZN(_02735_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06292_ (.A1(_02637_),
    .A2(_02733_),
    .B(_02735_),
    .ZN(_00137_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06293_ (.A1(\u_cpu.rf_ram.memory[1][2] ),
    .A2(_02733_),
    .ZN(_02736_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06294_ (.A1(_02642_),
    .A2(_02733_),
    .B(_02736_),
    .ZN(_00138_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06295_ (.A1(\u_cpu.rf_ram.memory[1][3] ),
    .A2(_02733_),
    .ZN(_02737_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06296_ (.A1(_02647_),
    .A2(_02733_),
    .B(_02737_),
    .ZN(_00139_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06297_ (.A1(\u_cpu.rf_ram.memory[1][4] ),
    .A2(_02733_),
    .ZN(_02738_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06298_ (.A1(_02652_),
    .A2(_02733_),
    .B(_02738_),
    .ZN(_00140_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06299_ (.A1(\u_cpu.rf_ram.memory[1][5] ),
    .A2(_02733_),
    .ZN(_02739_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06300_ (.A1(_02657_),
    .A2(_02733_),
    .B(_02739_),
    .ZN(_00141_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06301_ (.A1(\u_cpu.rf_ram.memory[1][6] ),
    .A2(_02733_),
    .ZN(_02740_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06302_ (.A1(_02662_),
    .A2(_02733_),
    .B(_02740_),
    .ZN(_00142_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06303_ (.A1(\u_cpu.rf_ram.memory[1][7] ),
    .A2(_02733_),
    .ZN(_02741_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06304_ (.A1(_02667_),
    .A2(_02733_),
    .B(_02741_),
    .ZN(_00143_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06305_ (.A1(_02616_),
    .A2(_02671_),
    .ZN(_02742_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06306_ (.A1(_02674_),
    .A2(_02742_),
    .ZN(_02743_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06307_ (.A1(_02731_),
    .A2(_02743_),
    .ZN(_02744_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06308_ (.I(_02744_),
    .ZN(_02745_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06309_ (.A1(\u_cpu.rf_ram.memory[7][0] ),
    .A2(_02745_),
    .ZN(_02746_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06310_ (.A1(_02632_),
    .A2(_02745_),
    .B(_02746_),
    .ZN(_00144_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06311_ (.A1(\u_cpu.rf_ram.memory[7][1] ),
    .A2(_02745_),
    .ZN(_02747_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06312_ (.A1(_02637_),
    .A2(_02745_),
    .B(_02747_),
    .ZN(_00145_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06313_ (.A1(\u_cpu.rf_ram.memory[7][2] ),
    .A2(_02745_),
    .ZN(_02748_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06314_ (.A1(_02642_),
    .A2(_02745_),
    .B(_02748_),
    .ZN(_00146_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06315_ (.A1(\u_cpu.rf_ram.memory[7][3] ),
    .A2(_02745_),
    .ZN(_02749_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06316_ (.A1(_02647_),
    .A2(_02745_),
    .B(_02749_),
    .ZN(_00147_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06317_ (.A1(\u_cpu.rf_ram.memory[7][4] ),
    .A2(_02745_),
    .ZN(_02750_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06318_ (.A1(_02652_),
    .A2(_02745_),
    .B(_02750_),
    .ZN(_00148_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06319_ (.A1(\u_cpu.rf_ram.memory[7][5] ),
    .A2(_02745_),
    .ZN(_02751_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06320_ (.A1(_02657_),
    .A2(_02745_),
    .B(_02751_),
    .ZN(_00149_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06321_ (.A1(\u_cpu.rf_ram.memory[7][6] ),
    .A2(_02745_),
    .ZN(_02752_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06322_ (.A1(_02662_),
    .A2(_02745_),
    .B(_02752_),
    .ZN(_00150_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06323_ (.A1(\u_cpu.rf_ram.memory[7][7] ),
    .A2(_02745_),
    .ZN(_02753_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06324_ (.A1(_02667_),
    .A2(_02745_),
    .B(_02753_),
    .ZN(_00151_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06325_ (.A1(_02614_),
    .A2(_02716_),
    .ZN(_02754_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06326_ (.A1(_02626_),
    .A2(_02754_),
    .ZN(_02755_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06327_ (.I(_02755_),
    .Z(_02756_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06328_ (.A1(\u_cpu.rf_ram.memory[80][0] ),
    .A2(_02756_),
    .ZN(_02757_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06329_ (.A1(_02669_),
    .A2(_02756_),
    .B(_02757_),
    .ZN(_00152_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06330_ (.A1(\u_cpu.rf_ram.memory[80][1] ),
    .A2(_02756_),
    .ZN(_02758_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06331_ (.A1(_02681_),
    .A2(_02756_),
    .B(_02758_),
    .ZN(_00153_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06332_ (.A1(\u_cpu.rf_ram.memory[80][2] ),
    .A2(_02756_),
    .ZN(_02759_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06333_ (.A1(_02683_),
    .A2(_02756_),
    .B(_02759_),
    .ZN(_00154_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06334_ (.A1(\u_cpu.rf_ram.memory[80][3] ),
    .A2(_02756_),
    .ZN(_02760_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06335_ (.A1(_02685_),
    .A2(_02756_),
    .B(_02760_),
    .ZN(_00155_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06336_ (.A1(\u_cpu.rf_ram.memory[80][4] ),
    .A2(_02756_),
    .ZN(_02761_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06337_ (.A1(_02687_),
    .A2(_02756_),
    .B(_02761_),
    .ZN(_00156_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06338_ (.A1(\u_cpu.rf_ram.memory[80][5] ),
    .A2(_02756_),
    .ZN(_02762_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06339_ (.A1(_02689_),
    .A2(_02756_),
    .B(_02762_),
    .ZN(_00157_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06340_ (.A1(\u_cpu.rf_ram.memory[80][6] ),
    .A2(_02756_),
    .ZN(_02763_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06341_ (.A1(_02691_),
    .A2(_02756_),
    .B(_02763_),
    .ZN(_00158_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06342_ (.A1(\u_cpu.rf_ram.memory[80][7] ),
    .A2(_02756_),
    .ZN(_02764_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06343_ (.A1(_02693_),
    .A2(_02756_),
    .B(_02764_),
    .ZN(_00159_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06344_ (.A1(_02609_),
    .A2(_02613_),
    .ZN(_02765_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06345_ (.A1(_02618_),
    .A2(_02765_),
    .ZN(_02766_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _06346_ (.A1(_02728_),
    .A2(_02608_),
    .A3(_02623_),
    .A4(_02729_),
    .Z(_02767_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06347_ (.I(_02767_),
    .Z(_02768_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06348_ (.A1(_02766_),
    .A2(_02768_),
    .ZN(_02769_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06349_ (.I(_02769_),
    .Z(_02770_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06350_ (.A1(\u_cpu.rf_ram.memory[78][0] ),
    .A2(_02770_),
    .ZN(_02771_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06351_ (.A1(_02669_),
    .A2(_02770_),
    .B(_02771_),
    .ZN(_00160_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06352_ (.A1(\u_cpu.rf_ram.memory[78][1] ),
    .A2(_02770_),
    .ZN(_02772_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06353_ (.A1(_02681_),
    .A2(_02770_),
    .B(_02772_),
    .ZN(_00161_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06354_ (.A1(\u_cpu.rf_ram.memory[78][2] ),
    .A2(_02770_),
    .ZN(_02773_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06355_ (.A1(_02683_),
    .A2(_02770_),
    .B(_02773_),
    .ZN(_00162_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06356_ (.A1(\u_cpu.rf_ram.memory[78][3] ),
    .A2(_02770_),
    .ZN(_02774_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06357_ (.A1(_02685_),
    .A2(_02770_),
    .B(_02774_),
    .ZN(_00163_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06358_ (.A1(\u_cpu.rf_ram.memory[78][4] ),
    .A2(_02770_),
    .ZN(_02775_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06359_ (.A1(_02687_),
    .A2(_02770_),
    .B(_02775_),
    .ZN(_00164_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06360_ (.A1(\u_cpu.rf_ram.memory[78][5] ),
    .A2(_02770_),
    .ZN(_02776_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06361_ (.A1(_02689_),
    .A2(_02770_),
    .B(_02776_),
    .ZN(_00165_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06362_ (.A1(\u_cpu.rf_ram.memory[78][6] ),
    .A2(_02770_),
    .ZN(_02777_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06363_ (.A1(_02691_),
    .A2(_02770_),
    .B(_02777_),
    .ZN(_00166_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06364_ (.A1(\u_cpu.rf_ram.memory[78][7] ),
    .A2(_02770_),
    .ZN(_02778_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06365_ (.A1(_02693_),
    .A2(_02770_),
    .B(_02778_),
    .ZN(_00167_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _06366_ (.A1(_02609_),
    .A2(_02673_),
    .Z(_02779_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06367_ (.A1(_02618_),
    .A2(_02779_),
    .ZN(_02780_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _06368_ (.A1(\u_cpu.cpu.immdec.imm11_7[2] ),
    .A2(\u_cpu.cpu.immdec.imm11_7[4] ),
    .A3(_02622_),
    .A4(_02729_),
    .ZN(_02781_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06369_ (.I(_02781_),
    .Z(_02782_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06370_ (.A1(_02780_),
    .A2(_02782_),
    .ZN(_02783_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06371_ (.I(_02783_),
    .Z(_02784_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06372_ (.A1(\u_cpu.rf_ram.memory[42][0] ),
    .A2(_02784_),
    .ZN(_02785_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06373_ (.A1(_02669_),
    .A2(_02784_),
    .B(_02785_),
    .ZN(_00168_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06374_ (.A1(\u_cpu.rf_ram.memory[42][1] ),
    .A2(_02784_),
    .ZN(_02786_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06375_ (.A1(_02681_),
    .A2(_02784_),
    .B(_02786_),
    .ZN(_00169_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06376_ (.A1(\u_cpu.rf_ram.memory[42][2] ),
    .A2(_02784_),
    .ZN(_02787_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06377_ (.A1(_02683_),
    .A2(_02784_),
    .B(_02787_),
    .ZN(_00170_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06378_ (.A1(\u_cpu.rf_ram.memory[42][3] ),
    .A2(_02784_),
    .ZN(_02788_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06379_ (.A1(_02685_),
    .A2(_02784_),
    .B(_02788_),
    .ZN(_00171_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06380_ (.A1(\u_cpu.rf_ram.memory[42][4] ),
    .A2(_02784_),
    .ZN(_02789_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06381_ (.A1(_02687_),
    .A2(_02784_),
    .B(_02789_),
    .ZN(_00172_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06382_ (.A1(\u_cpu.rf_ram.memory[42][5] ),
    .A2(_02784_),
    .ZN(_02790_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06383_ (.A1(_02689_),
    .A2(_02784_),
    .B(_02790_),
    .ZN(_00173_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06384_ (.A1(\u_cpu.rf_ram.memory[42][6] ),
    .A2(_02784_),
    .ZN(_02791_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06385_ (.A1(_02691_),
    .A2(_02784_),
    .B(_02791_),
    .ZN(_00174_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06386_ (.A1(\u_cpu.rf_ram.memory[42][7] ),
    .A2(_02784_),
    .ZN(_02792_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06387_ (.A1(_02693_),
    .A2(_02784_),
    .B(_02792_),
    .ZN(_00175_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06388_ (.A1(_02766_),
    .A2(_02782_),
    .ZN(_02793_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06389_ (.I(_02793_),
    .Z(_02794_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06390_ (.A1(\u_cpu.rf_ram.memory[46][0] ),
    .A2(_02794_),
    .ZN(_02795_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06391_ (.A1(_02669_),
    .A2(_02794_),
    .B(_02795_),
    .ZN(_00176_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06392_ (.A1(\u_cpu.rf_ram.memory[46][1] ),
    .A2(_02794_),
    .ZN(_02796_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06393_ (.A1(_02681_),
    .A2(_02794_),
    .B(_02796_),
    .ZN(_00177_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06394_ (.A1(\u_cpu.rf_ram.memory[46][2] ),
    .A2(_02794_),
    .ZN(_02797_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06395_ (.A1(_02683_),
    .A2(_02794_),
    .B(_02797_),
    .ZN(_00178_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06396_ (.A1(\u_cpu.rf_ram.memory[46][3] ),
    .A2(_02794_),
    .ZN(_02798_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06397_ (.A1(_02685_),
    .A2(_02794_),
    .B(_02798_),
    .ZN(_00179_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06398_ (.A1(\u_cpu.rf_ram.memory[46][4] ),
    .A2(_02794_),
    .ZN(_02799_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06399_ (.A1(_02687_),
    .A2(_02794_),
    .B(_02799_),
    .ZN(_00180_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06400_ (.A1(\u_cpu.rf_ram.memory[46][5] ),
    .A2(_02794_),
    .ZN(_02800_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06401_ (.A1(_02689_),
    .A2(_02794_),
    .B(_02800_),
    .ZN(_00181_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06402_ (.A1(\u_cpu.rf_ram.memory[46][6] ),
    .A2(_02794_),
    .ZN(_02801_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06403_ (.A1(_02691_),
    .A2(_02794_),
    .B(_02801_),
    .ZN(_00182_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06404_ (.A1(\u_cpu.rf_ram.memory[46][7] ),
    .A2(_02794_),
    .ZN(_02802_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06405_ (.A1(_02693_),
    .A2(_02794_),
    .B(_02802_),
    .ZN(_00183_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06406_ (.A1(_02672_),
    .A2(_02765_),
    .ZN(_02803_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06407_ (.A1(_02782_),
    .A2(_02803_),
    .ZN(_02804_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06408_ (.I(_02804_),
    .Z(_02805_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06409_ (.A1(\u_cpu.rf_ram.memory[45][0] ),
    .A2(_02805_),
    .ZN(_02806_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06410_ (.A1(_02669_),
    .A2(_02805_),
    .B(_02806_),
    .ZN(_00184_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06411_ (.A1(\u_cpu.rf_ram.memory[45][1] ),
    .A2(_02805_),
    .ZN(_02807_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06412_ (.A1(_02681_),
    .A2(_02805_),
    .B(_02807_),
    .ZN(_00185_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06413_ (.A1(\u_cpu.rf_ram.memory[45][2] ),
    .A2(_02805_),
    .ZN(_02808_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06414_ (.A1(_02683_),
    .A2(_02805_),
    .B(_02808_),
    .ZN(_00186_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06415_ (.A1(\u_cpu.rf_ram.memory[45][3] ),
    .A2(_02805_),
    .ZN(_02809_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06416_ (.A1(_02685_),
    .A2(_02805_),
    .B(_02809_),
    .ZN(_00187_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06417_ (.A1(\u_cpu.rf_ram.memory[45][4] ),
    .A2(_02805_),
    .ZN(_02810_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06418_ (.A1(_02687_),
    .A2(_02805_),
    .B(_02810_),
    .ZN(_00188_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06419_ (.A1(\u_cpu.rf_ram.memory[45][5] ),
    .A2(_02805_),
    .ZN(_02811_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06420_ (.A1(_02689_),
    .A2(_02805_),
    .B(_02811_),
    .ZN(_00189_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06421_ (.A1(\u_cpu.rf_ram.memory[45][6] ),
    .A2(_02805_),
    .ZN(_02812_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06422_ (.A1(_02691_),
    .A2(_02805_),
    .B(_02812_),
    .ZN(_00190_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06423_ (.A1(\u_cpu.rf_ram.memory[45][7] ),
    .A2(_02805_),
    .ZN(_02813_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06424_ (.A1(_02693_),
    .A2(_02805_),
    .B(_02813_),
    .ZN(_00191_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06425_ (.A1(_02716_),
    .A2(_02765_),
    .ZN(_02814_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06426_ (.A1(_02782_),
    .A2(_02814_),
    .ZN(_02815_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06427_ (.I(_02815_),
    .Z(_02816_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06428_ (.A1(\u_cpu.rf_ram.memory[44][0] ),
    .A2(_02816_),
    .ZN(_02817_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06429_ (.A1(_02669_),
    .A2(_02816_),
    .B(_02817_),
    .ZN(_00192_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06430_ (.A1(\u_cpu.rf_ram.memory[44][1] ),
    .A2(_02816_),
    .ZN(_02818_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06431_ (.A1(_02681_),
    .A2(_02816_),
    .B(_02818_),
    .ZN(_00193_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06432_ (.A1(\u_cpu.rf_ram.memory[44][2] ),
    .A2(_02816_),
    .ZN(_02819_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06433_ (.A1(_02683_),
    .A2(_02816_),
    .B(_02819_),
    .ZN(_00194_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06434_ (.A1(\u_cpu.rf_ram.memory[44][3] ),
    .A2(_02816_),
    .ZN(_02820_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06435_ (.A1(_02685_),
    .A2(_02816_),
    .B(_02820_),
    .ZN(_00195_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06436_ (.A1(\u_cpu.rf_ram.memory[44][4] ),
    .A2(_02816_),
    .ZN(_02821_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06437_ (.A1(_02687_),
    .A2(_02816_),
    .B(_02821_),
    .ZN(_00196_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06438_ (.A1(\u_cpu.rf_ram.memory[44][5] ),
    .A2(_02816_),
    .ZN(_02822_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06439_ (.A1(_02689_),
    .A2(_02816_),
    .B(_02822_),
    .ZN(_00197_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06440_ (.A1(\u_cpu.rf_ram.memory[44][6] ),
    .A2(_02816_),
    .ZN(_02823_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06441_ (.A1(_02691_),
    .A2(_02816_),
    .B(_02823_),
    .ZN(_00198_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06442_ (.A1(\u_cpu.rf_ram.memory[44][7] ),
    .A2(_02816_),
    .ZN(_02824_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06443_ (.A1(_02693_),
    .A2(_02816_),
    .B(_02824_),
    .ZN(_00199_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06444_ (.A1(_02614_),
    .A2(_02742_),
    .ZN(_02825_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _06445_ (.A1(_02728_),
    .A2(\u_cpu.cpu.immdec.imm11_7[4] ),
    .A3(_02622_),
    .A4(_02729_),
    .ZN(_02826_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06446_ (.I(_02826_),
    .Z(_02827_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06447_ (.A1(_02825_),
    .A2(_02827_),
    .ZN(_02828_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06448_ (.I(_02828_),
    .Z(_02829_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06449_ (.A1(\u_cpu.rf_ram.memory[51][0] ),
    .A2(_02829_),
    .ZN(_02830_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06450_ (.A1(_02669_),
    .A2(_02829_),
    .B(_02830_),
    .ZN(_00200_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06451_ (.A1(\u_cpu.rf_ram.memory[51][1] ),
    .A2(_02829_),
    .ZN(_02831_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06452_ (.A1(_02681_),
    .A2(_02829_),
    .B(_02831_),
    .ZN(_00201_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06453_ (.A1(\u_cpu.rf_ram.memory[51][2] ),
    .A2(_02829_),
    .ZN(_02832_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06454_ (.A1(_02683_),
    .A2(_02829_),
    .B(_02832_),
    .ZN(_00202_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06455_ (.A1(\u_cpu.rf_ram.memory[51][3] ),
    .A2(_02829_),
    .ZN(_02833_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06456_ (.A1(_02685_),
    .A2(_02829_),
    .B(_02833_),
    .ZN(_00203_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06457_ (.A1(\u_cpu.rf_ram.memory[51][4] ),
    .A2(_02829_),
    .ZN(_02834_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06458_ (.A1(_02687_),
    .A2(_02829_),
    .B(_02834_),
    .ZN(_00204_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06459_ (.A1(\u_cpu.rf_ram.memory[51][5] ),
    .A2(_02829_),
    .ZN(_02835_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06460_ (.A1(_02689_),
    .A2(_02829_),
    .B(_02835_),
    .ZN(_00205_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06461_ (.A1(\u_cpu.rf_ram.memory[51][6] ),
    .A2(_02829_),
    .ZN(_02836_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06462_ (.A1(_02691_),
    .A2(_02829_),
    .B(_02836_),
    .ZN(_00206_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06463_ (.A1(\u_cpu.rf_ram.memory[51][7] ),
    .A2(_02829_),
    .ZN(_02837_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06464_ (.A1(_02693_),
    .A2(_02829_),
    .B(_02837_),
    .ZN(_00207_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06465_ (.A1(_02672_),
    .A2(_02779_),
    .ZN(_02838_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06466_ (.A1(_02782_),
    .A2(_02838_),
    .ZN(_02839_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06467_ (.I(_02839_),
    .Z(_02840_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06468_ (.A1(\u_cpu.rf_ram.memory[41][0] ),
    .A2(_02840_),
    .ZN(_02841_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06469_ (.A1(_02669_),
    .A2(_02840_),
    .B(_02841_),
    .ZN(_00208_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06470_ (.A1(\u_cpu.rf_ram.memory[41][1] ),
    .A2(_02840_),
    .ZN(_02842_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06471_ (.A1(_02681_),
    .A2(_02840_),
    .B(_02842_),
    .ZN(_00209_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06472_ (.A1(\u_cpu.rf_ram.memory[41][2] ),
    .A2(_02840_),
    .ZN(_02843_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06473_ (.A1(_02683_),
    .A2(_02840_),
    .B(_02843_),
    .ZN(_00210_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06474_ (.A1(\u_cpu.rf_ram.memory[41][3] ),
    .A2(_02840_),
    .ZN(_02844_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06475_ (.A1(_02685_),
    .A2(_02840_),
    .B(_02844_),
    .ZN(_00211_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06476_ (.A1(\u_cpu.rf_ram.memory[41][4] ),
    .A2(_02840_),
    .ZN(_02845_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06477_ (.A1(_02687_),
    .A2(_02840_),
    .B(_02845_),
    .ZN(_00212_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06478_ (.A1(\u_cpu.rf_ram.memory[41][5] ),
    .A2(_02840_),
    .ZN(_02846_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06479_ (.A1(_02689_),
    .A2(_02840_),
    .B(_02846_),
    .ZN(_00213_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06480_ (.A1(\u_cpu.rf_ram.memory[41][6] ),
    .A2(_02840_),
    .ZN(_02847_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06481_ (.A1(_02691_),
    .A2(_02840_),
    .B(_02847_),
    .ZN(_00214_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06482_ (.A1(\u_cpu.rf_ram.memory[41][7] ),
    .A2(_02840_),
    .ZN(_02848_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06483_ (.A1(_02693_),
    .A2(_02840_),
    .B(_02848_),
    .ZN(_00215_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06484_ (.A1(_02742_),
    .A2(_02779_),
    .ZN(_02849_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06485_ (.A1(_02782_),
    .A2(_02849_),
    .ZN(_02850_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06486_ (.I(_02850_),
    .Z(_02851_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06487_ (.A1(\u_cpu.rf_ram.memory[43][0] ),
    .A2(_02851_),
    .ZN(_02852_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06488_ (.A1(_02669_),
    .A2(_02851_),
    .B(_02852_),
    .ZN(_00216_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06489_ (.A1(\u_cpu.rf_ram.memory[43][1] ),
    .A2(_02851_),
    .ZN(_02853_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06490_ (.A1(_02681_),
    .A2(_02851_),
    .B(_02853_),
    .ZN(_00217_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06491_ (.A1(\u_cpu.rf_ram.memory[43][2] ),
    .A2(_02851_),
    .ZN(_02854_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06492_ (.A1(_02683_),
    .A2(_02851_),
    .B(_02854_),
    .ZN(_00218_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06493_ (.A1(\u_cpu.rf_ram.memory[43][3] ),
    .A2(_02851_),
    .ZN(_02855_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06494_ (.A1(_02685_),
    .A2(_02851_),
    .B(_02855_),
    .ZN(_00219_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06495_ (.A1(\u_cpu.rf_ram.memory[43][4] ),
    .A2(_02851_),
    .ZN(_02856_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06496_ (.A1(_02687_),
    .A2(_02851_),
    .B(_02856_),
    .ZN(_00220_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06497_ (.A1(\u_cpu.rf_ram.memory[43][5] ),
    .A2(_02851_),
    .ZN(_02857_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06498_ (.A1(_02689_),
    .A2(_02851_),
    .B(_02857_),
    .ZN(_00221_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06499_ (.A1(\u_cpu.rf_ram.memory[43][6] ),
    .A2(_02851_),
    .ZN(_02858_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06500_ (.A1(_02691_),
    .A2(_02851_),
    .B(_02858_),
    .ZN(_00222_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06501_ (.A1(\u_cpu.rf_ram.memory[43][7] ),
    .A2(_02851_),
    .ZN(_02859_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06502_ (.A1(_02693_),
    .A2(_02851_),
    .B(_02859_),
    .ZN(_00223_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06503_ (.A1(_02754_),
    .A2(_02827_),
    .ZN(_02860_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06504_ (.I(_02860_),
    .Z(_02861_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06505_ (.A1(\u_cpu.rf_ram.memory[48][0] ),
    .A2(_02861_),
    .ZN(_02862_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06506_ (.A1(_02669_),
    .A2(_02861_),
    .B(_02862_),
    .ZN(_00224_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06507_ (.A1(\u_cpu.rf_ram.memory[48][1] ),
    .A2(_02861_),
    .ZN(_02863_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06508_ (.A1(_02681_),
    .A2(_02861_),
    .B(_02863_),
    .ZN(_00225_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06509_ (.A1(\u_cpu.rf_ram.memory[48][2] ),
    .A2(_02861_),
    .ZN(_02864_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06510_ (.A1(_02683_),
    .A2(_02861_),
    .B(_02864_),
    .ZN(_00226_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06511_ (.A1(\u_cpu.rf_ram.memory[48][3] ),
    .A2(_02861_),
    .ZN(_02865_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06512_ (.A1(_02685_),
    .A2(_02861_),
    .B(_02865_),
    .ZN(_00227_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06513_ (.A1(\u_cpu.rf_ram.memory[48][4] ),
    .A2(_02861_),
    .ZN(_02866_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06514_ (.A1(_02687_),
    .A2(_02861_),
    .B(_02866_),
    .ZN(_00228_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06515_ (.A1(\u_cpu.rf_ram.memory[48][5] ),
    .A2(_02861_),
    .ZN(_02867_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06516_ (.A1(_02689_),
    .A2(_02861_),
    .B(_02867_),
    .ZN(_00229_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06517_ (.A1(\u_cpu.rf_ram.memory[48][6] ),
    .A2(_02861_),
    .ZN(_02868_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06518_ (.A1(_02691_),
    .A2(_02861_),
    .B(_02868_),
    .ZN(_00230_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06519_ (.A1(\u_cpu.rf_ram.memory[48][7] ),
    .A2(_02861_),
    .ZN(_02869_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06520_ (.A1(_02693_),
    .A2(_02861_),
    .B(_02869_),
    .ZN(_00231_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06521_ (.A1(_02742_),
    .A2(_02765_),
    .ZN(_02870_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06522_ (.A1(_02782_),
    .A2(_02870_),
    .ZN(_02871_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06523_ (.I(_02871_),
    .Z(_02872_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06524_ (.A1(\u_cpu.rf_ram.memory[47][0] ),
    .A2(_02872_),
    .ZN(_02873_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06525_ (.A1(_02669_),
    .A2(_02872_),
    .B(_02873_),
    .ZN(_00232_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06526_ (.A1(\u_cpu.rf_ram.memory[47][1] ),
    .A2(_02872_),
    .ZN(_02874_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06527_ (.A1(_02681_),
    .A2(_02872_),
    .B(_02874_),
    .ZN(_00233_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06528_ (.A1(\u_cpu.rf_ram.memory[47][2] ),
    .A2(_02872_),
    .ZN(_02875_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06529_ (.A1(_02683_),
    .A2(_02872_),
    .B(_02875_),
    .ZN(_00234_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06530_ (.A1(\u_cpu.rf_ram.memory[47][3] ),
    .A2(_02872_),
    .ZN(_02876_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06531_ (.A1(_02685_),
    .A2(_02872_),
    .B(_02876_),
    .ZN(_00235_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06532_ (.A1(\u_cpu.rf_ram.memory[47][4] ),
    .A2(_02872_),
    .ZN(_02877_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06533_ (.A1(_02687_),
    .A2(_02872_),
    .B(_02877_),
    .ZN(_00236_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06534_ (.A1(\u_cpu.rf_ram.memory[47][5] ),
    .A2(_02872_),
    .ZN(_02878_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06535_ (.A1(_02689_),
    .A2(_02872_),
    .B(_02878_),
    .ZN(_00237_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06536_ (.A1(\u_cpu.rf_ram.memory[47][6] ),
    .A2(_02872_),
    .ZN(_02879_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06537_ (.A1(_02691_),
    .A2(_02872_),
    .B(_02879_),
    .ZN(_00238_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06538_ (.A1(\u_cpu.rf_ram.memory[47][7] ),
    .A2(_02872_),
    .ZN(_02880_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06539_ (.A1(_02693_),
    .A2(_02872_),
    .B(_02880_),
    .ZN(_00239_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06540_ (.I(_02631_),
    .Z(_02881_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06541_ (.A1(_02619_),
    .A2(_02827_),
    .ZN(_02882_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06542_ (.I(_02882_),
    .Z(_02883_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06543_ (.A1(\u_cpu.rf_ram.memory[50][0] ),
    .A2(_02883_),
    .ZN(_02884_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06544_ (.A1(_02881_),
    .A2(_02883_),
    .B(_02884_),
    .ZN(_00240_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06545_ (.I(_02636_),
    .Z(_02885_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06546_ (.A1(\u_cpu.rf_ram.memory[50][1] ),
    .A2(_02883_),
    .ZN(_02886_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06547_ (.A1(_02885_),
    .A2(_02883_),
    .B(_02886_),
    .ZN(_00241_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06548_ (.I(_02641_),
    .Z(_02887_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06549_ (.A1(\u_cpu.rf_ram.memory[50][2] ),
    .A2(_02883_),
    .ZN(_02888_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06550_ (.A1(_02887_),
    .A2(_02883_),
    .B(_02888_),
    .ZN(_00242_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06551_ (.I(_02646_),
    .Z(_02889_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06552_ (.A1(\u_cpu.rf_ram.memory[50][3] ),
    .A2(_02883_),
    .ZN(_02890_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06553_ (.A1(_02889_),
    .A2(_02883_),
    .B(_02890_),
    .ZN(_00243_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06554_ (.I(_02651_),
    .Z(_02891_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06555_ (.A1(\u_cpu.rf_ram.memory[50][4] ),
    .A2(_02883_),
    .ZN(_02892_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06556_ (.A1(_02891_),
    .A2(_02883_),
    .B(_02892_),
    .ZN(_00244_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06557_ (.I(_02656_),
    .Z(_02893_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06558_ (.A1(\u_cpu.rf_ram.memory[50][5] ),
    .A2(_02883_),
    .ZN(_02894_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06559_ (.A1(_02893_),
    .A2(_02883_),
    .B(_02894_),
    .ZN(_00245_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06560_ (.I(_02661_),
    .Z(_02895_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06561_ (.A1(\u_cpu.rf_ram.memory[50][6] ),
    .A2(_02883_),
    .ZN(_02896_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06562_ (.A1(_02895_),
    .A2(_02883_),
    .B(_02896_),
    .ZN(_00246_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06563_ (.I(_02666_),
    .Z(_02897_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06564_ (.A1(\u_cpu.rf_ram.memory[50][7] ),
    .A2(_02883_),
    .ZN(_02898_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06565_ (.A1(_02897_),
    .A2(_02883_),
    .B(_02898_),
    .ZN(_00247_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06566_ (.A1(_02717_),
    .A2(_02731_),
    .ZN(_02899_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06567_ (.I(_02899_),
    .ZN(_02900_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06568_ (.A1(\u_cpu.rf_ram.memory[4][0] ),
    .A2(_02900_),
    .ZN(_02901_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06569_ (.A1(_02632_),
    .A2(_02900_),
    .B(_02901_),
    .ZN(_00248_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06570_ (.A1(\u_cpu.rf_ram.memory[4][1] ),
    .A2(_02900_),
    .ZN(_02902_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06571_ (.A1(_02637_),
    .A2(_02900_),
    .B(_02902_),
    .ZN(_00249_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06572_ (.A1(\u_cpu.rf_ram.memory[4][2] ),
    .A2(_02900_),
    .ZN(_02903_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06573_ (.A1(_02642_),
    .A2(_02900_),
    .B(_02903_),
    .ZN(_00250_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06574_ (.A1(\u_cpu.rf_ram.memory[4][3] ),
    .A2(_02900_),
    .ZN(_02904_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06575_ (.A1(_02647_),
    .A2(_02900_),
    .B(_02904_),
    .ZN(_00251_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06576_ (.A1(\u_cpu.rf_ram.memory[4][4] ),
    .A2(_02900_),
    .ZN(_02905_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06577_ (.A1(_02652_),
    .A2(_02900_),
    .B(_02905_),
    .ZN(_00252_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06578_ (.A1(\u_cpu.rf_ram.memory[4][5] ),
    .A2(_02900_),
    .ZN(_02906_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06579_ (.A1(_02657_),
    .A2(_02900_),
    .B(_02906_),
    .ZN(_00253_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06580_ (.A1(\u_cpu.rf_ram.memory[4][6] ),
    .A2(_02900_),
    .ZN(_02907_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06581_ (.A1(_02662_),
    .A2(_02900_),
    .B(_02907_),
    .ZN(_00254_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06582_ (.A1(\u_cpu.rf_ram.memory[4][7] ),
    .A2(_02900_),
    .ZN(_02908_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06583_ (.A1(_02667_),
    .A2(_02900_),
    .B(_02908_),
    .ZN(_00255_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _06584_ (.I(_02464_),
    .ZN(_02909_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06585_ (.A1(\u_arbiter.i_wb_cpu_ack ),
    .A2(_02461_),
    .ZN(_02910_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06586_ (.A1(_02909_),
    .A2(\u_arbiter.i_wb_cpu_ibus_adr[1] ),
    .B(_02910_),
    .ZN(_02911_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06587_ (.A1(\u_cpu.cpu.state.genblk1.misalign_trap_sync_r ),
    .A2(\u_cpu.cpu.state.stage_two_req ),
    .B(_02911_),
    .ZN(_02912_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06588_ (.A1(_02395_),
    .A2(_02912_),
    .ZN(_00256_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06589_ (.A1(_01444_),
    .A2(_02285_),
    .ZN(_02913_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06590_ (.A1(_02307_),
    .A2(_02311_),
    .Z(_02914_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06591_ (.A1(_02913_),
    .A2(_02914_),
    .ZN(_02915_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _06592_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[3] ),
    .A2(\u_arbiter.i_wb_cpu_dbus_dat[2] ),
    .A3(\u_arbiter.i_wb_cpu_dbus_dat[0] ),
    .A4(\u_arbiter.i_wb_cpu_dbus_dat[1] ),
    .Z(_02916_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06593_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[4] ),
    .A2(_02916_),
    .ZN(_02917_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06594_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[5] ),
    .A2(_02917_),
    .Z(_02918_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06595_ (.A1(_02915_),
    .A2(_02918_),
    .ZN(_02919_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06596_ (.A1(_02263_),
    .A2(_02598_),
    .B(_02314_),
    .ZN(_02920_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06597_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[6] ),
    .A2(_02920_),
    .ZN(_02921_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06598_ (.A1(_02919_),
    .A2(_02921_),
    .ZN(_02922_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _06599_ (.A1(_01441_),
    .A2(_02309_),
    .A3(_02922_),
    .ZN(_02923_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06600_ (.A1(\u_arbiter.i_wb_cpu_ack ),
    .A2(_02397_),
    .ZN(_02924_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06601_ (.A1(_02313_),
    .A2(_02923_),
    .B(_02924_),
    .ZN(_02925_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06602_ (.A1(\u_cpu.cpu.state.genblk1.misalign_trap_sync_r ),
    .A2(_02393_),
    .ZN(_02926_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06603_ (.A1(_02305_),
    .A2(_02925_),
    .B(_02926_),
    .ZN(_02927_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06604_ (.A1(_02912_),
    .A2(_02927_),
    .ZN(_02928_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06605_ (.A1(\u_cpu.rf_ram_if.rcnt[0] ),
    .A2(_02928_),
    .ZN(_00257_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _06606_ (.A1(\u_cpu.rf_ram_if.rcnt[0] ),
    .A2(\u_cpu.rf_ram_if.rcnt[2] ),
    .A3(\u_cpu.rf_ram_if.rcnt[1] ),
    .Z(_02929_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _06607_ (.A1(_02615_),
    .A2(_02928_),
    .A3(_02929_),
    .ZN(_00258_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06608_ (.A1(_01634_),
    .A2(_02929_),
    .ZN(_02930_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _06609_ (.A1(_01634_),
    .A2(_02929_),
    .Z(_02931_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _06610_ (.A1(_02912_),
    .A2(_02927_),
    .A3(_02930_),
    .A4(_02931_),
    .Z(_02932_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06611_ (.I(_02932_),
    .Z(_00259_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06612_ (.A1(_01635_),
    .A2(_02930_),
    .Z(_02933_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06613_ (.A1(_02928_),
    .A2(_02933_),
    .ZN(_00260_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06614_ (.A1(_02677_),
    .A2(_02754_),
    .ZN(_02934_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06615_ (.I(_02934_),
    .Z(_02935_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06616_ (.A1(\u_cpu.rf_ram.memory[16][0] ),
    .A2(_02935_),
    .ZN(_02936_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06617_ (.A1(_02881_),
    .A2(_02935_),
    .B(_02936_),
    .ZN(_00261_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06618_ (.A1(\u_cpu.rf_ram.memory[16][1] ),
    .A2(_02935_),
    .ZN(_02937_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06619_ (.A1(_02885_),
    .A2(_02935_),
    .B(_02937_),
    .ZN(_00262_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06620_ (.A1(\u_cpu.rf_ram.memory[16][2] ),
    .A2(_02935_),
    .ZN(_02938_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06621_ (.A1(_02887_),
    .A2(_02935_),
    .B(_02938_),
    .ZN(_00263_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06622_ (.A1(\u_cpu.rf_ram.memory[16][3] ),
    .A2(_02935_),
    .ZN(_02939_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06623_ (.A1(_02889_),
    .A2(_02935_),
    .B(_02939_),
    .ZN(_00264_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06624_ (.A1(\u_cpu.rf_ram.memory[16][4] ),
    .A2(_02935_),
    .ZN(_02940_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06625_ (.A1(_02891_),
    .A2(_02935_),
    .B(_02940_),
    .ZN(_00265_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06626_ (.A1(\u_cpu.rf_ram.memory[16][5] ),
    .A2(_02935_),
    .ZN(_02941_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06627_ (.A1(_02893_),
    .A2(_02935_),
    .B(_02941_),
    .ZN(_00266_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06628_ (.A1(\u_cpu.rf_ram.memory[16][6] ),
    .A2(_02935_),
    .ZN(_02942_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06629_ (.A1(_02895_),
    .A2(_02935_),
    .B(_02942_),
    .ZN(_00267_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06630_ (.A1(\u_cpu.rf_ram.memory[16][7] ),
    .A2(_02935_),
    .ZN(_02943_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06631_ (.A1(_02897_),
    .A2(_02935_),
    .B(_02943_),
    .ZN(_00268_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06632_ (.A1(_02677_),
    .A2(_02695_),
    .ZN(_02944_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06633_ (.I(_02944_),
    .Z(_02945_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06634_ (.A1(\u_cpu.rf_ram.memory[17][0] ),
    .A2(_02945_),
    .ZN(_02946_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06635_ (.A1(_02881_),
    .A2(_02945_),
    .B(_02946_),
    .ZN(_00269_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06636_ (.A1(\u_cpu.rf_ram.memory[17][1] ),
    .A2(_02945_),
    .ZN(_02947_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06637_ (.A1(_02885_),
    .A2(_02945_),
    .B(_02947_),
    .ZN(_00270_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06638_ (.A1(\u_cpu.rf_ram.memory[17][2] ),
    .A2(_02945_),
    .ZN(_02948_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06639_ (.A1(_02887_),
    .A2(_02945_),
    .B(_02948_),
    .ZN(_00271_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06640_ (.A1(\u_cpu.rf_ram.memory[17][3] ),
    .A2(_02945_),
    .ZN(_02949_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06641_ (.A1(_02889_),
    .A2(_02945_),
    .B(_02949_),
    .ZN(_00272_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06642_ (.A1(\u_cpu.rf_ram.memory[17][4] ),
    .A2(_02945_),
    .ZN(_02950_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06643_ (.A1(_02891_),
    .A2(_02945_),
    .B(_02950_),
    .ZN(_00273_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06644_ (.A1(\u_cpu.rf_ram.memory[17][5] ),
    .A2(_02945_),
    .ZN(_02951_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06645_ (.A1(_02893_),
    .A2(_02945_),
    .B(_02951_),
    .ZN(_00274_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06646_ (.A1(\u_cpu.rf_ram.memory[17][6] ),
    .A2(_02945_),
    .ZN(_02952_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06647_ (.A1(_02895_),
    .A2(_02945_),
    .B(_02952_),
    .ZN(_00275_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06648_ (.A1(\u_cpu.rf_ram.memory[17][7] ),
    .A2(_02945_),
    .ZN(_02953_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06649_ (.A1(_02897_),
    .A2(_02945_),
    .B(_02953_),
    .ZN(_00276_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06650_ (.A1(_02716_),
    .A2(_02779_),
    .ZN(_02954_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06651_ (.A1(_02782_),
    .A2(_02954_),
    .ZN(_02955_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06652_ (.I(_02955_),
    .Z(_02956_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06653_ (.A1(\u_cpu.rf_ram.memory[40][0] ),
    .A2(_02956_),
    .ZN(_02957_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06654_ (.A1(_02881_),
    .A2(_02956_),
    .B(_02957_),
    .ZN(_00277_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06655_ (.A1(\u_cpu.rf_ram.memory[40][1] ),
    .A2(_02956_),
    .ZN(_02958_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06656_ (.A1(_02885_),
    .A2(_02956_),
    .B(_02958_),
    .ZN(_00278_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06657_ (.A1(\u_cpu.rf_ram.memory[40][2] ),
    .A2(_02956_),
    .ZN(_02959_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06658_ (.A1(_02887_),
    .A2(_02956_),
    .B(_02959_),
    .ZN(_00279_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06659_ (.A1(\u_cpu.rf_ram.memory[40][3] ),
    .A2(_02956_),
    .ZN(_02960_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06660_ (.A1(_02889_),
    .A2(_02956_),
    .B(_02960_),
    .ZN(_00280_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06661_ (.A1(\u_cpu.rf_ram.memory[40][4] ),
    .A2(_02956_),
    .ZN(_02961_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06662_ (.A1(_02891_),
    .A2(_02956_),
    .B(_02961_),
    .ZN(_00281_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06663_ (.A1(\u_cpu.rf_ram.memory[40][5] ),
    .A2(_02956_),
    .ZN(_02962_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06664_ (.A1(_02893_),
    .A2(_02956_),
    .B(_02962_),
    .ZN(_00282_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06665_ (.A1(\u_cpu.rf_ram.memory[40][6] ),
    .A2(_02956_),
    .ZN(_02963_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06666_ (.A1(_02895_),
    .A2(_02956_),
    .B(_02963_),
    .ZN(_00283_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06667_ (.A1(\u_cpu.rf_ram.memory[40][7] ),
    .A2(_02956_),
    .ZN(_02964_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06668_ (.A1(_02897_),
    .A2(_02956_),
    .B(_02964_),
    .ZN(_00284_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _06669_ (.A1(_02728_),
    .A2(_02624_),
    .A3(_02729_),
    .ZN(_02965_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06670_ (.A1(_02743_),
    .A2(_02965_),
    .ZN(_02966_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06671_ (.I(_02966_),
    .Z(_02967_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06672_ (.A1(\u_cpu.rf_ram.memory[119][0] ),
    .A2(_02967_),
    .ZN(_02968_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06673_ (.A1(_02881_),
    .A2(_02967_),
    .B(_02968_),
    .ZN(_00285_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06674_ (.A1(\u_cpu.rf_ram.memory[119][1] ),
    .A2(_02967_),
    .ZN(_02969_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06675_ (.A1(_02885_),
    .A2(_02967_),
    .B(_02969_),
    .ZN(_00286_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06676_ (.A1(\u_cpu.rf_ram.memory[119][2] ),
    .A2(_02967_),
    .ZN(_02970_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06677_ (.A1(_02887_),
    .A2(_02967_),
    .B(_02970_),
    .ZN(_00287_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06678_ (.A1(\u_cpu.rf_ram.memory[119][3] ),
    .A2(_02967_),
    .ZN(_02971_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06679_ (.A1(_02889_),
    .A2(_02967_),
    .B(_02971_),
    .ZN(_00288_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06680_ (.A1(\u_cpu.rf_ram.memory[119][4] ),
    .A2(_02967_),
    .ZN(_02972_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06681_ (.A1(_02891_),
    .A2(_02967_),
    .B(_02972_),
    .ZN(_00289_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06682_ (.A1(\u_cpu.rf_ram.memory[119][5] ),
    .A2(_02967_),
    .ZN(_02973_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06683_ (.A1(_02893_),
    .A2(_02967_),
    .B(_02973_),
    .ZN(_00290_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06684_ (.A1(\u_cpu.rf_ram.memory[119][6] ),
    .A2(_02967_),
    .ZN(_02974_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06685_ (.A1(_02895_),
    .A2(_02967_),
    .B(_02974_),
    .ZN(_00291_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06686_ (.A1(\u_cpu.rf_ram.memory[119][7] ),
    .A2(_02967_),
    .ZN(_02975_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06687_ (.A1(_02897_),
    .A2(_02967_),
    .B(_02975_),
    .ZN(_00292_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06688_ (.A1(_02608_),
    .A2(_02622_),
    .ZN(_02976_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06689_ (.A1(_02695_),
    .A2(_02976_),
    .ZN(_02977_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06690_ (.I(_02977_),
    .Z(_02978_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06691_ (.A1(\u_cpu.rf_ram.memory[129][0] ),
    .A2(_02978_),
    .ZN(_02979_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06692_ (.A1(_02881_),
    .A2(_02978_),
    .B(_02979_),
    .ZN(_00293_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06693_ (.A1(\u_cpu.rf_ram.memory[129][1] ),
    .A2(_02978_),
    .ZN(_02980_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06694_ (.A1(_02885_),
    .A2(_02978_),
    .B(_02980_),
    .ZN(_00294_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06695_ (.A1(\u_cpu.rf_ram.memory[129][2] ),
    .A2(_02978_),
    .ZN(_02981_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06696_ (.A1(_02887_),
    .A2(_02978_),
    .B(_02981_),
    .ZN(_00295_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06697_ (.A1(\u_cpu.rf_ram.memory[129][3] ),
    .A2(_02978_),
    .ZN(_02982_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06698_ (.A1(_02889_),
    .A2(_02978_),
    .B(_02982_),
    .ZN(_00296_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06699_ (.A1(\u_cpu.rf_ram.memory[129][4] ),
    .A2(_02978_),
    .ZN(_02983_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06700_ (.A1(_02891_),
    .A2(_02978_),
    .B(_02983_),
    .ZN(_00297_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06701_ (.A1(\u_cpu.rf_ram.memory[129][5] ),
    .A2(_02978_),
    .ZN(_02984_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06702_ (.A1(_02893_),
    .A2(_02978_),
    .B(_02984_),
    .ZN(_00298_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06703_ (.A1(\u_cpu.rf_ram.memory[129][6] ),
    .A2(_02978_),
    .ZN(_02985_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06704_ (.A1(_02895_),
    .A2(_02978_),
    .B(_02985_),
    .ZN(_00299_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06705_ (.A1(\u_cpu.rf_ram.memory[129][7] ),
    .A2(_02978_),
    .ZN(_02986_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06706_ (.A1(_02897_),
    .A2(_02978_),
    .B(_02986_),
    .ZN(_00300_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06707_ (.A1(_02849_),
    .A2(_02976_),
    .ZN(_02987_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06708_ (.I(_02987_),
    .Z(_02988_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06709_ (.A1(\u_cpu.rf_ram.memory[139][0] ),
    .A2(_02988_),
    .ZN(_02989_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06710_ (.A1(_02881_),
    .A2(_02988_),
    .B(_02989_),
    .ZN(_00301_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06711_ (.A1(\u_cpu.rf_ram.memory[139][1] ),
    .A2(_02988_),
    .ZN(_02990_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06712_ (.A1(_02885_),
    .A2(_02988_),
    .B(_02990_),
    .ZN(_00302_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06713_ (.A1(\u_cpu.rf_ram.memory[139][2] ),
    .A2(_02988_),
    .ZN(_02991_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06714_ (.A1(_02887_),
    .A2(_02988_),
    .B(_02991_),
    .ZN(_00303_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06715_ (.A1(\u_cpu.rf_ram.memory[139][3] ),
    .A2(_02988_),
    .ZN(_02992_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06716_ (.A1(_02889_),
    .A2(_02988_),
    .B(_02992_),
    .ZN(_00304_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06717_ (.A1(\u_cpu.rf_ram.memory[139][4] ),
    .A2(_02988_),
    .ZN(_02993_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06718_ (.A1(_02891_),
    .A2(_02988_),
    .B(_02993_),
    .ZN(_00305_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06719_ (.A1(\u_cpu.rf_ram.memory[139][5] ),
    .A2(_02988_),
    .ZN(_02994_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06720_ (.A1(_02893_),
    .A2(_02988_),
    .B(_02994_),
    .ZN(_00306_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06721_ (.A1(\u_cpu.rf_ram.memory[139][6] ),
    .A2(_02988_),
    .ZN(_02995_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06722_ (.A1(_02895_),
    .A2(_02988_),
    .B(_02995_),
    .ZN(_00307_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06723_ (.A1(\u_cpu.rf_ram.memory[139][7] ),
    .A2(_02988_),
    .ZN(_02996_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06724_ (.A1(_02897_),
    .A2(_02988_),
    .B(_02996_),
    .ZN(_00308_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06725_ (.A1(_02768_),
    .A2(_02803_),
    .ZN(_02997_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06726_ (.I(_02997_),
    .Z(_02998_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06727_ (.A1(\u_cpu.rf_ram.memory[77][0] ),
    .A2(_02998_),
    .ZN(_02999_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06728_ (.A1(_02881_),
    .A2(_02998_),
    .B(_02999_),
    .ZN(_00309_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06729_ (.A1(\u_cpu.rf_ram.memory[77][1] ),
    .A2(_02998_),
    .ZN(_03000_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06730_ (.A1(_02885_),
    .A2(_02998_),
    .B(_03000_),
    .ZN(_00310_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06731_ (.A1(\u_cpu.rf_ram.memory[77][2] ),
    .A2(_02998_),
    .ZN(_03001_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06732_ (.A1(_02887_),
    .A2(_02998_),
    .B(_03001_),
    .ZN(_00311_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06733_ (.A1(\u_cpu.rf_ram.memory[77][3] ),
    .A2(_02998_),
    .ZN(_03002_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06734_ (.A1(_02889_),
    .A2(_02998_),
    .B(_03002_),
    .ZN(_00312_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06735_ (.A1(\u_cpu.rf_ram.memory[77][4] ),
    .A2(_02998_),
    .ZN(_03003_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06736_ (.A1(_02891_),
    .A2(_02998_),
    .B(_03003_),
    .ZN(_00313_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06737_ (.A1(\u_cpu.rf_ram.memory[77][5] ),
    .A2(_02998_),
    .ZN(_03004_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06738_ (.A1(_02893_),
    .A2(_02998_),
    .B(_03004_),
    .ZN(_00314_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06739_ (.A1(\u_cpu.rf_ram.memory[77][6] ),
    .A2(_02998_),
    .ZN(_03005_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06740_ (.A1(_02895_),
    .A2(_02998_),
    .B(_03005_),
    .ZN(_00315_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06741_ (.A1(\u_cpu.rf_ram.memory[77][7] ),
    .A2(_02998_),
    .ZN(_03006_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06742_ (.A1(_02897_),
    .A2(_02998_),
    .B(_03006_),
    .ZN(_00316_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06743_ (.A1(_02768_),
    .A2(_02780_),
    .ZN(_03007_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06744_ (.I(_03007_),
    .Z(_03008_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06745_ (.A1(\u_cpu.rf_ram.memory[74][0] ),
    .A2(_03008_),
    .ZN(_03009_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06746_ (.A1(_02881_),
    .A2(_03008_),
    .B(_03009_),
    .ZN(_00317_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06747_ (.A1(\u_cpu.rf_ram.memory[74][1] ),
    .A2(_03008_),
    .ZN(_03010_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06748_ (.A1(_02885_),
    .A2(_03008_),
    .B(_03010_),
    .ZN(_00318_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06749_ (.A1(\u_cpu.rf_ram.memory[74][2] ),
    .A2(_03008_),
    .ZN(_03011_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06750_ (.A1(_02887_),
    .A2(_03008_),
    .B(_03011_),
    .ZN(_00319_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06751_ (.A1(\u_cpu.rf_ram.memory[74][3] ),
    .A2(_03008_),
    .ZN(_03012_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06752_ (.A1(_02889_),
    .A2(_03008_),
    .B(_03012_),
    .ZN(_00320_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06753_ (.A1(\u_cpu.rf_ram.memory[74][4] ),
    .A2(_03008_),
    .ZN(_03013_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06754_ (.A1(_02891_),
    .A2(_03008_),
    .B(_03013_),
    .ZN(_00321_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06755_ (.A1(\u_cpu.rf_ram.memory[74][5] ),
    .A2(_03008_),
    .ZN(_03014_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06756_ (.A1(_02893_),
    .A2(_03008_),
    .B(_03014_),
    .ZN(_00322_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06757_ (.A1(\u_cpu.rf_ram.memory[74][6] ),
    .A2(_03008_),
    .ZN(_03015_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06758_ (.A1(_02895_),
    .A2(_03008_),
    .B(_03015_),
    .ZN(_00323_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06759_ (.A1(\u_cpu.rf_ram.memory[74][7] ),
    .A2(_03008_),
    .ZN(_03016_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06760_ (.A1(_02897_),
    .A2(_03008_),
    .B(_03016_),
    .ZN(_00324_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06761_ (.A1(_02768_),
    .A2(_02814_),
    .ZN(_03017_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06762_ (.I(_03017_),
    .Z(_03018_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06763_ (.A1(\u_cpu.rf_ram.memory[76][0] ),
    .A2(_03018_),
    .ZN(_03019_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06764_ (.A1(_02881_),
    .A2(_03018_),
    .B(_03019_),
    .ZN(_00325_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06765_ (.A1(\u_cpu.rf_ram.memory[76][1] ),
    .A2(_03018_),
    .ZN(_03020_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06766_ (.A1(_02885_),
    .A2(_03018_),
    .B(_03020_),
    .ZN(_00326_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06767_ (.A1(\u_cpu.rf_ram.memory[76][2] ),
    .A2(_03018_),
    .ZN(_03021_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06768_ (.A1(_02887_),
    .A2(_03018_),
    .B(_03021_),
    .ZN(_00327_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06769_ (.A1(\u_cpu.rf_ram.memory[76][3] ),
    .A2(_03018_),
    .ZN(_03022_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06770_ (.A1(_02889_),
    .A2(_03018_),
    .B(_03022_),
    .ZN(_00328_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06771_ (.A1(\u_cpu.rf_ram.memory[76][4] ),
    .A2(_03018_),
    .ZN(_03023_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06772_ (.A1(_02891_),
    .A2(_03018_),
    .B(_03023_),
    .ZN(_00329_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06773_ (.A1(\u_cpu.rf_ram.memory[76][5] ),
    .A2(_03018_),
    .ZN(_03024_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06774_ (.A1(_02893_),
    .A2(_03018_),
    .B(_03024_),
    .ZN(_00330_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06775_ (.A1(\u_cpu.rf_ram.memory[76][6] ),
    .A2(_03018_),
    .ZN(_03025_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06776_ (.A1(_02895_),
    .A2(_03018_),
    .B(_03025_),
    .ZN(_00331_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06777_ (.A1(\u_cpu.rf_ram.memory[76][7] ),
    .A2(_03018_),
    .ZN(_03026_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06778_ (.A1(_02897_),
    .A2(_03018_),
    .B(_03026_),
    .ZN(_00332_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06779_ (.A1(_02768_),
    .A2(_02849_),
    .ZN(_03027_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06780_ (.I(_03027_),
    .Z(_03028_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06781_ (.A1(\u_cpu.rf_ram.memory[75][0] ),
    .A2(_03028_),
    .ZN(_03029_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06782_ (.A1(_02881_),
    .A2(_03028_),
    .B(_03029_),
    .ZN(_00333_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06783_ (.A1(\u_cpu.rf_ram.memory[75][1] ),
    .A2(_03028_),
    .ZN(_03030_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06784_ (.A1(_02885_),
    .A2(_03028_),
    .B(_03030_),
    .ZN(_00334_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06785_ (.A1(\u_cpu.rf_ram.memory[75][2] ),
    .A2(_03028_),
    .ZN(_03031_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06786_ (.A1(_02887_),
    .A2(_03028_),
    .B(_03031_),
    .ZN(_00335_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06787_ (.A1(\u_cpu.rf_ram.memory[75][3] ),
    .A2(_03028_),
    .ZN(_03032_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06788_ (.A1(_02889_),
    .A2(_03028_),
    .B(_03032_),
    .ZN(_00336_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06789_ (.A1(\u_cpu.rf_ram.memory[75][4] ),
    .A2(_03028_),
    .ZN(_03033_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06790_ (.A1(_02891_),
    .A2(_03028_),
    .B(_03033_),
    .ZN(_00337_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06791_ (.A1(\u_cpu.rf_ram.memory[75][5] ),
    .A2(_03028_),
    .ZN(_03034_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06792_ (.A1(_02893_),
    .A2(_03028_),
    .B(_03034_),
    .ZN(_00338_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06793_ (.A1(\u_cpu.rf_ram.memory[75][6] ),
    .A2(_03028_),
    .ZN(_03035_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06794_ (.A1(_02895_),
    .A2(_03028_),
    .B(_03035_),
    .ZN(_00339_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06795_ (.A1(\u_cpu.rf_ram.memory[75][7] ),
    .A2(_03028_),
    .ZN(_03036_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06796_ (.A1(_02897_),
    .A2(_03028_),
    .B(_03036_),
    .ZN(_00340_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06797_ (.A1(_02618_),
    .A2(_02674_),
    .ZN(_03037_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06798_ (.A1(_02731_),
    .A2(_03037_),
    .ZN(_03038_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06799_ (.I(_03038_),
    .ZN(_03039_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06800_ (.A1(\u_cpu.rf_ram.memory[6][0] ),
    .A2(_03039_),
    .ZN(_03040_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06801_ (.A1(_02632_),
    .A2(_03039_),
    .B(_03040_),
    .ZN(_00341_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06802_ (.A1(\u_cpu.rf_ram.memory[6][1] ),
    .A2(_03039_),
    .ZN(_03041_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06803_ (.A1(_02637_),
    .A2(_03039_),
    .B(_03041_),
    .ZN(_00342_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06804_ (.A1(\u_cpu.rf_ram.memory[6][2] ),
    .A2(_03039_),
    .ZN(_03042_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06805_ (.A1(_02642_),
    .A2(_03039_),
    .B(_03042_),
    .ZN(_00343_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06806_ (.A1(\u_cpu.rf_ram.memory[6][3] ),
    .A2(_03039_),
    .ZN(_03043_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06807_ (.A1(_02647_),
    .A2(_03039_),
    .B(_03043_),
    .ZN(_00344_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06808_ (.A1(\u_cpu.rf_ram.memory[6][4] ),
    .A2(_03039_),
    .ZN(_03044_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06809_ (.A1(_02652_),
    .A2(_03039_),
    .B(_03044_),
    .ZN(_00345_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06810_ (.A1(\u_cpu.rf_ram.memory[6][5] ),
    .A2(_03039_),
    .ZN(_03045_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06811_ (.A1(_02657_),
    .A2(_03039_),
    .B(_03045_),
    .ZN(_00346_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06812_ (.A1(\u_cpu.rf_ram.memory[6][6] ),
    .A2(_03039_),
    .ZN(_03046_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06813_ (.A1(_02662_),
    .A2(_03039_),
    .B(_03046_),
    .ZN(_00347_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06814_ (.A1(\u_cpu.rf_ram.memory[6][7] ),
    .A2(_03039_),
    .ZN(_03047_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06815_ (.A1(_02667_),
    .A2(_03039_),
    .B(_03047_),
    .ZN(_00348_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06816_ (.A1(_02717_),
    .A2(_02768_),
    .ZN(_03048_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06817_ (.I(_03048_),
    .Z(_03049_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06818_ (.A1(\u_cpu.rf_ram.memory[68][0] ),
    .A2(_03049_),
    .ZN(_03050_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06819_ (.A1(_02881_),
    .A2(_03049_),
    .B(_03050_),
    .ZN(_00349_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06820_ (.A1(\u_cpu.rf_ram.memory[68][1] ),
    .A2(_03049_),
    .ZN(_03051_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06821_ (.A1(_02885_),
    .A2(_03049_),
    .B(_03051_),
    .ZN(_00350_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06822_ (.A1(\u_cpu.rf_ram.memory[68][2] ),
    .A2(_03049_),
    .ZN(_03052_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06823_ (.A1(_02887_),
    .A2(_03049_),
    .B(_03052_),
    .ZN(_00351_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06824_ (.A1(\u_cpu.rf_ram.memory[68][3] ),
    .A2(_03049_),
    .ZN(_03053_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06825_ (.A1(_02889_),
    .A2(_03049_),
    .B(_03053_),
    .ZN(_00352_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06826_ (.A1(\u_cpu.rf_ram.memory[68][4] ),
    .A2(_03049_),
    .ZN(_03054_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06827_ (.A1(_02891_),
    .A2(_03049_),
    .B(_03054_),
    .ZN(_00353_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06828_ (.A1(\u_cpu.rf_ram.memory[68][5] ),
    .A2(_03049_),
    .ZN(_03055_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06829_ (.A1(_02893_),
    .A2(_03049_),
    .B(_03055_),
    .ZN(_00354_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06830_ (.A1(\u_cpu.rf_ram.memory[68][6] ),
    .A2(_03049_),
    .ZN(_03056_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06831_ (.A1(_02895_),
    .A2(_03049_),
    .B(_03056_),
    .ZN(_00355_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06832_ (.A1(\u_cpu.rf_ram.memory[68][7] ),
    .A2(_03049_),
    .ZN(_03057_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06833_ (.A1(_02897_),
    .A2(_03049_),
    .B(_03057_),
    .ZN(_00356_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06834_ (.A1(_02768_),
    .A2(_02825_),
    .ZN(_03058_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06835_ (.I(_03058_),
    .Z(_03059_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06836_ (.A1(\u_cpu.rf_ram.memory[67][0] ),
    .A2(_03059_),
    .ZN(_03060_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06837_ (.A1(_02881_),
    .A2(_03059_),
    .B(_03060_),
    .ZN(_00357_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06838_ (.A1(\u_cpu.rf_ram.memory[67][1] ),
    .A2(_03059_),
    .ZN(_03061_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06839_ (.A1(_02885_),
    .A2(_03059_),
    .B(_03061_),
    .ZN(_00358_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06840_ (.A1(\u_cpu.rf_ram.memory[67][2] ),
    .A2(_03059_),
    .ZN(_03062_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06841_ (.A1(_02887_),
    .A2(_03059_),
    .B(_03062_),
    .ZN(_00359_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06842_ (.A1(\u_cpu.rf_ram.memory[67][3] ),
    .A2(_03059_),
    .ZN(_03063_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06843_ (.A1(_02889_),
    .A2(_03059_),
    .B(_03063_),
    .ZN(_00360_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06844_ (.A1(\u_cpu.rf_ram.memory[67][4] ),
    .A2(_03059_),
    .ZN(_03064_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06845_ (.A1(_02891_),
    .A2(_03059_),
    .B(_03064_),
    .ZN(_00361_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06846_ (.A1(\u_cpu.rf_ram.memory[67][5] ),
    .A2(_03059_),
    .ZN(_03065_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06847_ (.A1(_02893_),
    .A2(_03059_),
    .B(_03065_),
    .ZN(_00362_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06848_ (.A1(\u_cpu.rf_ram.memory[67][6] ),
    .A2(_03059_),
    .ZN(_03066_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06849_ (.A1(_02895_),
    .A2(_03059_),
    .B(_03066_),
    .ZN(_00363_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06850_ (.A1(\u_cpu.rf_ram.memory[67][7] ),
    .A2(_03059_),
    .ZN(_03067_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06851_ (.A1(_02897_),
    .A2(_03059_),
    .B(_03067_),
    .ZN(_00364_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06852_ (.A1(_02619_),
    .A2(_02768_),
    .ZN(_03068_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06853_ (.I(_03068_),
    .Z(_03069_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06854_ (.A1(\u_cpu.rf_ram.memory[66][0] ),
    .A2(_03069_),
    .ZN(_03070_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06855_ (.A1(_02881_),
    .A2(_03069_),
    .B(_03070_),
    .ZN(_00365_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06856_ (.A1(\u_cpu.rf_ram.memory[66][1] ),
    .A2(_03069_),
    .ZN(_03071_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06857_ (.A1(_02885_),
    .A2(_03069_),
    .B(_03071_),
    .ZN(_00366_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06858_ (.A1(\u_cpu.rf_ram.memory[66][2] ),
    .A2(_03069_),
    .ZN(_03072_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06859_ (.A1(_02887_),
    .A2(_03069_),
    .B(_03072_),
    .ZN(_00367_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06860_ (.A1(\u_cpu.rf_ram.memory[66][3] ),
    .A2(_03069_),
    .ZN(_03073_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06861_ (.A1(_02889_),
    .A2(_03069_),
    .B(_03073_),
    .ZN(_00368_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06862_ (.A1(\u_cpu.rf_ram.memory[66][4] ),
    .A2(_03069_),
    .ZN(_03074_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06863_ (.A1(_02891_),
    .A2(_03069_),
    .B(_03074_),
    .ZN(_00369_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06864_ (.A1(\u_cpu.rf_ram.memory[66][5] ),
    .A2(_03069_),
    .ZN(_03075_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06865_ (.A1(_02893_),
    .A2(_03069_),
    .B(_03075_),
    .ZN(_00370_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06866_ (.A1(\u_cpu.rf_ram.memory[66][6] ),
    .A2(_03069_),
    .ZN(_03076_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06867_ (.A1(_02895_),
    .A2(_03069_),
    .B(_03076_),
    .ZN(_00371_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06868_ (.A1(\u_cpu.rf_ram.memory[66][7] ),
    .A2(_03069_),
    .ZN(_03077_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06869_ (.A1(_02897_),
    .A2(_03069_),
    .B(_03077_),
    .ZN(_00372_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06870_ (.A1(_02695_),
    .A2(_02768_),
    .ZN(_03078_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06871_ (.I(_03078_),
    .Z(_03079_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06872_ (.A1(\u_cpu.rf_ram.memory[65][0] ),
    .A2(_03079_),
    .ZN(_03080_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06873_ (.A1(_02881_),
    .A2(_03079_),
    .B(_03080_),
    .ZN(_00373_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06874_ (.A1(\u_cpu.rf_ram.memory[65][1] ),
    .A2(_03079_),
    .ZN(_03081_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06875_ (.A1(_02885_),
    .A2(_03079_),
    .B(_03081_),
    .ZN(_00374_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06876_ (.A1(\u_cpu.rf_ram.memory[65][2] ),
    .A2(_03079_),
    .ZN(_03082_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06877_ (.A1(_02887_),
    .A2(_03079_),
    .B(_03082_),
    .ZN(_00375_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06878_ (.A1(\u_cpu.rf_ram.memory[65][3] ),
    .A2(_03079_),
    .ZN(_03083_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06879_ (.A1(_02889_),
    .A2(_03079_),
    .B(_03083_),
    .ZN(_00376_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06880_ (.A1(\u_cpu.rf_ram.memory[65][4] ),
    .A2(_03079_),
    .ZN(_03084_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06881_ (.A1(_02891_),
    .A2(_03079_),
    .B(_03084_),
    .ZN(_00377_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06882_ (.A1(\u_cpu.rf_ram.memory[65][5] ),
    .A2(_03079_),
    .ZN(_03085_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06883_ (.A1(_02893_),
    .A2(_03079_),
    .B(_03085_),
    .ZN(_00378_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06884_ (.A1(\u_cpu.rf_ram.memory[65][6] ),
    .A2(_03079_),
    .ZN(_03086_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06885_ (.A1(_02895_),
    .A2(_03079_),
    .B(_03086_),
    .ZN(_00379_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06886_ (.A1(\u_cpu.rf_ram.memory[65][7] ),
    .A2(_03079_),
    .ZN(_03087_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06887_ (.A1(_02897_),
    .A2(_03079_),
    .B(_03087_),
    .ZN(_00380_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06888_ (.A1(_02754_),
    .A2(_02768_),
    .ZN(_03088_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06889_ (.I(_03088_),
    .Z(_03089_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06890_ (.A1(\u_cpu.rf_ram.memory[64][0] ),
    .A2(_03089_),
    .ZN(_03090_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06891_ (.A1(_02881_),
    .A2(_03089_),
    .B(_03090_),
    .ZN(_00381_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06892_ (.A1(\u_cpu.rf_ram.memory[64][1] ),
    .A2(_03089_),
    .ZN(_03091_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06893_ (.A1(_02885_),
    .A2(_03089_),
    .B(_03091_),
    .ZN(_00382_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06894_ (.A1(\u_cpu.rf_ram.memory[64][2] ),
    .A2(_03089_),
    .ZN(_03092_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06895_ (.A1(_02887_),
    .A2(_03089_),
    .B(_03092_),
    .ZN(_00383_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06896_ (.A1(\u_cpu.rf_ram.memory[64][3] ),
    .A2(_03089_),
    .ZN(_03093_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06897_ (.A1(_02889_),
    .A2(_03089_),
    .B(_03093_),
    .ZN(_00384_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06898_ (.A1(\u_cpu.rf_ram.memory[64][4] ),
    .A2(_03089_),
    .ZN(_03094_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06899_ (.A1(_02891_),
    .A2(_03089_),
    .B(_03094_),
    .ZN(_00385_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06900_ (.A1(\u_cpu.rf_ram.memory[64][5] ),
    .A2(_03089_),
    .ZN(_03095_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06901_ (.A1(_02893_),
    .A2(_03089_),
    .B(_03095_),
    .ZN(_00386_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06902_ (.A1(\u_cpu.rf_ram.memory[64][6] ),
    .A2(_03089_),
    .ZN(_03096_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06903_ (.A1(_02895_),
    .A2(_03089_),
    .B(_03096_),
    .ZN(_00387_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06904_ (.A1(\u_cpu.rf_ram.memory[64][7] ),
    .A2(_03089_),
    .ZN(_03097_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06905_ (.A1(_02897_),
    .A2(_03089_),
    .B(_03097_),
    .ZN(_00388_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06906_ (.I(_02631_),
    .Z(_03098_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06907_ (.A1(_02677_),
    .A2(_02803_),
    .ZN(_03099_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06908_ (.I(_03099_),
    .Z(_03100_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06909_ (.A1(\u_cpu.rf_ram.memory[29][0] ),
    .A2(_03100_),
    .ZN(_03101_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06910_ (.A1(_03098_),
    .A2(_03100_),
    .B(_03101_),
    .ZN(_00389_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06911_ (.I(_02636_),
    .Z(_03102_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06912_ (.A1(\u_cpu.rf_ram.memory[29][1] ),
    .A2(_03100_),
    .ZN(_03103_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06913_ (.A1(_03102_),
    .A2(_03100_),
    .B(_03103_),
    .ZN(_00390_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06914_ (.I(_02641_),
    .Z(_03104_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06915_ (.A1(\u_cpu.rf_ram.memory[29][2] ),
    .A2(_03100_),
    .ZN(_03105_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06916_ (.A1(_03104_),
    .A2(_03100_),
    .B(_03105_),
    .ZN(_00391_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06917_ (.I(_02646_),
    .Z(_03106_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06918_ (.A1(\u_cpu.rf_ram.memory[29][3] ),
    .A2(_03100_),
    .ZN(_03107_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06919_ (.A1(_03106_),
    .A2(_03100_),
    .B(_03107_),
    .ZN(_00392_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06920_ (.I(_02651_),
    .Z(_03108_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06921_ (.A1(\u_cpu.rf_ram.memory[29][4] ),
    .A2(_03100_),
    .ZN(_03109_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06922_ (.A1(_03108_),
    .A2(_03100_),
    .B(_03109_),
    .ZN(_00393_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06923_ (.I(_02656_),
    .Z(_03110_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06924_ (.A1(\u_cpu.rf_ram.memory[29][5] ),
    .A2(_03100_),
    .ZN(_03111_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06925_ (.A1(_03110_),
    .A2(_03100_),
    .B(_03111_),
    .ZN(_00394_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06926_ (.I(_02661_),
    .Z(_03112_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06927_ (.A1(\u_cpu.rf_ram.memory[29][6] ),
    .A2(_03100_),
    .ZN(_03113_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06928_ (.A1(_03112_),
    .A2(_03100_),
    .B(_03113_),
    .ZN(_00395_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06929_ (.I(_02666_),
    .Z(_03114_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06930_ (.A1(\u_cpu.rf_ram.memory[29][7] ),
    .A2(_03100_),
    .ZN(_03115_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06931_ (.A1(_03114_),
    .A2(_03100_),
    .B(_03115_),
    .ZN(_00396_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06932_ (.A1(_02827_),
    .A2(_02870_),
    .ZN(_03116_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06933_ (.I(_03116_),
    .Z(_03117_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06934_ (.A1(\u_cpu.rf_ram.memory[63][0] ),
    .A2(_03117_),
    .ZN(_03118_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06935_ (.A1(_03098_),
    .A2(_03117_),
    .B(_03118_),
    .ZN(_00397_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06936_ (.A1(\u_cpu.rf_ram.memory[63][1] ),
    .A2(_03117_),
    .ZN(_03119_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06937_ (.A1(_03102_),
    .A2(_03117_),
    .B(_03119_),
    .ZN(_00398_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06938_ (.A1(\u_cpu.rf_ram.memory[63][2] ),
    .A2(_03117_),
    .ZN(_03120_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06939_ (.A1(_03104_),
    .A2(_03117_),
    .B(_03120_),
    .ZN(_00399_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06940_ (.A1(\u_cpu.rf_ram.memory[63][3] ),
    .A2(_03117_),
    .ZN(_03121_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06941_ (.A1(_03106_),
    .A2(_03117_),
    .B(_03121_),
    .ZN(_00400_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06942_ (.A1(\u_cpu.rf_ram.memory[63][4] ),
    .A2(_03117_),
    .ZN(_03122_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06943_ (.A1(_03108_),
    .A2(_03117_),
    .B(_03122_),
    .ZN(_00401_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06944_ (.A1(\u_cpu.rf_ram.memory[63][5] ),
    .A2(_03117_),
    .ZN(_03123_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06945_ (.A1(_03110_),
    .A2(_03117_),
    .B(_03123_),
    .ZN(_00402_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06946_ (.A1(\u_cpu.rf_ram.memory[63][6] ),
    .A2(_03117_),
    .ZN(_03124_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06947_ (.A1(_03112_),
    .A2(_03117_),
    .B(_03124_),
    .ZN(_00403_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06948_ (.A1(\u_cpu.rf_ram.memory[63][7] ),
    .A2(_03117_),
    .ZN(_03125_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06949_ (.A1(_03114_),
    .A2(_03117_),
    .B(_03125_),
    .ZN(_00404_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06950_ (.A1(_02766_),
    .A2(_02827_),
    .ZN(_03126_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06951_ (.I(_03126_),
    .Z(_03127_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06952_ (.A1(\u_cpu.rf_ram.memory[62][0] ),
    .A2(_03127_),
    .ZN(_03128_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06953_ (.A1(_03098_),
    .A2(_03127_),
    .B(_03128_),
    .ZN(_00405_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06954_ (.A1(\u_cpu.rf_ram.memory[62][1] ),
    .A2(_03127_),
    .ZN(_03129_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06955_ (.A1(_03102_),
    .A2(_03127_),
    .B(_03129_),
    .ZN(_00406_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06956_ (.A1(\u_cpu.rf_ram.memory[62][2] ),
    .A2(_03127_),
    .ZN(_03130_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06957_ (.A1(_03104_),
    .A2(_03127_),
    .B(_03130_),
    .ZN(_00407_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06958_ (.A1(\u_cpu.rf_ram.memory[62][3] ),
    .A2(_03127_),
    .ZN(_03131_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06959_ (.A1(_03106_),
    .A2(_03127_),
    .B(_03131_),
    .ZN(_00408_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06960_ (.A1(\u_cpu.rf_ram.memory[62][4] ),
    .A2(_03127_),
    .ZN(_03132_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06961_ (.A1(_03108_),
    .A2(_03127_),
    .B(_03132_),
    .ZN(_00409_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06962_ (.A1(\u_cpu.rf_ram.memory[62][5] ),
    .A2(_03127_),
    .ZN(_03133_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06963_ (.A1(_03110_),
    .A2(_03127_),
    .B(_03133_),
    .ZN(_00410_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06964_ (.A1(\u_cpu.rf_ram.memory[62][6] ),
    .A2(_03127_),
    .ZN(_03134_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06965_ (.A1(_03112_),
    .A2(_03127_),
    .B(_03134_),
    .ZN(_00411_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06966_ (.A1(\u_cpu.rf_ram.memory[62][7] ),
    .A2(_03127_),
    .ZN(_03135_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06967_ (.A1(_03114_),
    .A2(_03127_),
    .B(_03135_),
    .ZN(_00412_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06968_ (.A1(_02803_),
    .A2(_02827_),
    .ZN(_03136_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06969_ (.I(_03136_),
    .Z(_03137_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06970_ (.A1(\u_cpu.rf_ram.memory[61][0] ),
    .A2(_03137_),
    .ZN(_03138_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06971_ (.A1(_03098_),
    .A2(_03137_),
    .B(_03138_),
    .ZN(_00413_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06972_ (.A1(\u_cpu.rf_ram.memory[61][1] ),
    .A2(_03137_),
    .ZN(_03139_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06973_ (.A1(_03102_),
    .A2(_03137_),
    .B(_03139_),
    .ZN(_00414_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06974_ (.A1(\u_cpu.rf_ram.memory[61][2] ),
    .A2(_03137_),
    .ZN(_03140_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06975_ (.A1(_03104_),
    .A2(_03137_),
    .B(_03140_),
    .ZN(_00415_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06976_ (.A1(\u_cpu.rf_ram.memory[61][3] ),
    .A2(_03137_),
    .ZN(_03141_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06977_ (.A1(_03106_),
    .A2(_03137_),
    .B(_03141_),
    .ZN(_00416_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06978_ (.A1(\u_cpu.rf_ram.memory[61][4] ),
    .A2(_03137_),
    .ZN(_03142_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06979_ (.A1(_03108_),
    .A2(_03137_),
    .B(_03142_),
    .ZN(_00417_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06980_ (.A1(\u_cpu.rf_ram.memory[61][5] ),
    .A2(_03137_),
    .ZN(_03143_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06981_ (.A1(_03110_),
    .A2(_03137_),
    .B(_03143_),
    .ZN(_00418_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06982_ (.A1(\u_cpu.rf_ram.memory[61][6] ),
    .A2(_03137_),
    .ZN(_03144_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06983_ (.A1(_03112_),
    .A2(_03137_),
    .B(_03144_),
    .ZN(_00419_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06984_ (.A1(\u_cpu.rf_ram.memory[61][7] ),
    .A2(_03137_),
    .ZN(_03145_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06985_ (.A1(_03114_),
    .A2(_03137_),
    .B(_03145_),
    .ZN(_00420_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06986_ (.A1(_02814_),
    .A2(_02827_),
    .ZN(_03146_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06987_ (.I(_03146_),
    .Z(_03147_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06988_ (.A1(\u_cpu.rf_ram.memory[60][0] ),
    .A2(_03147_),
    .ZN(_03148_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06989_ (.A1(_03098_),
    .A2(_03147_),
    .B(_03148_),
    .ZN(_00421_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06990_ (.A1(\u_cpu.rf_ram.memory[60][1] ),
    .A2(_03147_),
    .ZN(_03149_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06991_ (.A1(_03102_),
    .A2(_03147_),
    .B(_03149_),
    .ZN(_00422_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06992_ (.A1(\u_cpu.rf_ram.memory[60][2] ),
    .A2(_03147_),
    .ZN(_03150_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06993_ (.A1(_03104_),
    .A2(_03147_),
    .B(_03150_),
    .ZN(_00423_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06994_ (.A1(\u_cpu.rf_ram.memory[60][3] ),
    .A2(_03147_),
    .ZN(_03151_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06995_ (.A1(_03106_),
    .A2(_03147_),
    .B(_03151_),
    .ZN(_00424_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06996_ (.A1(\u_cpu.rf_ram.memory[60][4] ),
    .A2(_03147_),
    .ZN(_03152_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06997_ (.A1(_03108_),
    .A2(_03147_),
    .B(_03152_),
    .ZN(_00425_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06998_ (.A1(\u_cpu.rf_ram.memory[60][5] ),
    .A2(_03147_),
    .ZN(_03153_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06999_ (.A1(_03110_),
    .A2(_03147_),
    .B(_03153_),
    .ZN(_00426_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07000_ (.A1(\u_cpu.rf_ram.memory[60][6] ),
    .A2(_03147_),
    .ZN(_03154_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07001_ (.A1(_03112_),
    .A2(_03147_),
    .B(_03154_),
    .ZN(_00427_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07002_ (.A1(\u_cpu.rf_ram.memory[60][7] ),
    .A2(_03147_),
    .ZN(_03155_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07003_ (.A1(_03114_),
    .A2(_03147_),
    .B(_03155_),
    .ZN(_00428_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07004_ (.A1(_02677_),
    .A2(_02825_),
    .ZN(_03156_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07005_ (.I(_03156_),
    .Z(_03157_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07006_ (.A1(\u_cpu.rf_ram.memory[19][0] ),
    .A2(_03157_),
    .ZN(_03158_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07007_ (.A1(_03098_),
    .A2(_03157_),
    .B(_03158_),
    .ZN(_00429_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07008_ (.A1(\u_cpu.rf_ram.memory[19][1] ),
    .A2(_03157_),
    .ZN(_03159_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07009_ (.A1(_03102_),
    .A2(_03157_),
    .B(_03159_),
    .ZN(_00430_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07010_ (.A1(\u_cpu.rf_ram.memory[19][2] ),
    .A2(_03157_),
    .ZN(_03160_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07011_ (.A1(_03104_),
    .A2(_03157_),
    .B(_03160_),
    .ZN(_00431_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07012_ (.A1(\u_cpu.rf_ram.memory[19][3] ),
    .A2(_03157_),
    .ZN(_03161_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07013_ (.A1(_03106_),
    .A2(_03157_),
    .B(_03161_),
    .ZN(_00432_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07014_ (.A1(\u_cpu.rf_ram.memory[19][4] ),
    .A2(_03157_),
    .ZN(_03162_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07015_ (.A1(_03108_),
    .A2(_03157_),
    .B(_03162_),
    .ZN(_00433_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07016_ (.A1(\u_cpu.rf_ram.memory[19][5] ),
    .A2(_03157_),
    .ZN(_03163_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07017_ (.A1(_03110_),
    .A2(_03157_),
    .B(_03163_),
    .ZN(_00434_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07018_ (.A1(\u_cpu.rf_ram.memory[19][6] ),
    .A2(_03157_),
    .ZN(_03164_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07019_ (.A1(_03112_),
    .A2(_03157_),
    .B(_03164_),
    .ZN(_00435_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07020_ (.A1(\u_cpu.rf_ram.memory[19][7] ),
    .A2(_03157_),
    .ZN(_03165_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07021_ (.A1(_03114_),
    .A2(_03157_),
    .B(_03165_),
    .ZN(_00436_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07022_ (.A1(_02675_),
    .A2(_02731_),
    .ZN(_03166_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07023_ (.I(_03166_),
    .ZN(_03167_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07024_ (.A1(\u_cpu.rf_ram.memory[5][0] ),
    .A2(_03167_),
    .ZN(_03168_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07025_ (.A1(_02632_),
    .A2(_03167_),
    .B(_03168_),
    .ZN(_00437_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07026_ (.A1(\u_cpu.rf_ram.memory[5][1] ),
    .A2(_03167_),
    .ZN(_03169_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07027_ (.A1(_02637_),
    .A2(_03167_),
    .B(_03169_),
    .ZN(_00438_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07028_ (.A1(\u_cpu.rf_ram.memory[5][2] ),
    .A2(_03167_),
    .ZN(_03170_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07029_ (.A1(_02642_),
    .A2(_03167_),
    .B(_03170_),
    .ZN(_00439_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07030_ (.A1(\u_cpu.rf_ram.memory[5][3] ),
    .A2(_03167_),
    .ZN(_03171_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07031_ (.A1(_02647_),
    .A2(_03167_),
    .B(_03171_),
    .ZN(_00440_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07032_ (.A1(\u_cpu.rf_ram.memory[5][4] ),
    .A2(_03167_),
    .ZN(_03172_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07033_ (.A1(_02652_),
    .A2(_03167_),
    .B(_03172_),
    .ZN(_00441_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07034_ (.A1(\u_cpu.rf_ram.memory[5][5] ),
    .A2(_03167_),
    .ZN(_03173_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07035_ (.A1(_02657_),
    .A2(_03167_),
    .B(_03173_),
    .ZN(_00442_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07036_ (.A1(\u_cpu.rf_ram.memory[5][6] ),
    .A2(_03167_),
    .ZN(_03174_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07037_ (.A1(_02662_),
    .A2(_03167_),
    .B(_03174_),
    .ZN(_00443_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07038_ (.A1(\u_cpu.rf_ram.memory[5][7] ),
    .A2(_03167_),
    .ZN(_03175_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07039_ (.A1(_02667_),
    .A2(_03167_),
    .B(_03175_),
    .ZN(_00444_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07040_ (.A1(_02780_),
    .A2(_02827_),
    .ZN(_03176_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07041_ (.I(_03176_),
    .Z(_03177_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07042_ (.A1(\u_cpu.rf_ram.memory[58][0] ),
    .A2(_03177_),
    .ZN(_03178_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07043_ (.A1(_03098_),
    .A2(_03177_),
    .B(_03178_),
    .ZN(_00445_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07044_ (.A1(\u_cpu.rf_ram.memory[58][1] ),
    .A2(_03177_),
    .ZN(_03179_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07045_ (.A1(_03102_),
    .A2(_03177_),
    .B(_03179_),
    .ZN(_00446_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07046_ (.A1(\u_cpu.rf_ram.memory[58][2] ),
    .A2(_03177_),
    .ZN(_03180_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07047_ (.A1(_03104_),
    .A2(_03177_),
    .B(_03180_),
    .ZN(_00447_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07048_ (.A1(\u_cpu.rf_ram.memory[58][3] ),
    .A2(_03177_),
    .ZN(_03181_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07049_ (.A1(_03106_),
    .A2(_03177_),
    .B(_03181_),
    .ZN(_00448_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07050_ (.A1(\u_cpu.rf_ram.memory[58][4] ),
    .A2(_03177_),
    .ZN(_03182_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07051_ (.A1(_03108_),
    .A2(_03177_),
    .B(_03182_),
    .ZN(_00449_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07052_ (.A1(\u_cpu.rf_ram.memory[58][5] ),
    .A2(_03177_),
    .ZN(_03183_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07053_ (.A1(_03110_),
    .A2(_03177_),
    .B(_03183_),
    .ZN(_00450_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07054_ (.A1(\u_cpu.rf_ram.memory[58][6] ),
    .A2(_03177_),
    .ZN(_03184_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07055_ (.A1(_03112_),
    .A2(_03177_),
    .B(_03184_),
    .ZN(_00451_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07056_ (.A1(\u_cpu.rf_ram.memory[58][7] ),
    .A2(_03177_),
    .ZN(_03185_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07057_ (.A1(_03114_),
    .A2(_03177_),
    .B(_03185_),
    .ZN(_00452_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07058_ (.A1(_02827_),
    .A2(_02838_),
    .ZN(_03186_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07059_ (.I(_03186_),
    .Z(_03187_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07060_ (.A1(\u_cpu.rf_ram.memory[57][0] ),
    .A2(_03187_),
    .ZN(_03188_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07061_ (.A1(_03098_),
    .A2(_03187_),
    .B(_03188_),
    .ZN(_00453_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07062_ (.A1(\u_cpu.rf_ram.memory[57][1] ),
    .A2(_03187_),
    .ZN(_03189_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07063_ (.A1(_03102_),
    .A2(_03187_),
    .B(_03189_),
    .ZN(_00454_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07064_ (.A1(\u_cpu.rf_ram.memory[57][2] ),
    .A2(_03187_),
    .ZN(_03190_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07065_ (.A1(_03104_),
    .A2(_03187_),
    .B(_03190_),
    .ZN(_00455_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07066_ (.A1(\u_cpu.rf_ram.memory[57][3] ),
    .A2(_03187_),
    .ZN(_03191_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07067_ (.A1(_03106_),
    .A2(_03187_),
    .B(_03191_),
    .ZN(_00456_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07068_ (.A1(\u_cpu.rf_ram.memory[57][4] ),
    .A2(_03187_),
    .ZN(_03192_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07069_ (.A1(_03108_),
    .A2(_03187_),
    .B(_03192_),
    .ZN(_00457_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07070_ (.A1(\u_cpu.rf_ram.memory[57][5] ),
    .A2(_03187_),
    .ZN(_03193_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07071_ (.A1(_03110_),
    .A2(_03187_),
    .B(_03193_),
    .ZN(_00458_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07072_ (.A1(\u_cpu.rf_ram.memory[57][6] ),
    .A2(_03187_),
    .ZN(_03194_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07073_ (.A1(_03112_),
    .A2(_03187_),
    .B(_03194_),
    .ZN(_00459_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07074_ (.A1(\u_cpu.rf_ram.memory[57][7] ),
    .A2(_03187_),
    .ZN(_03195_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07075_ (.A1(_03114_),
    .A2(_03187_),
    .B(_03195_),
    .ZN(_00460_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07076_ (.A1(_02827_),
    .A2(_02954_),
    .ZN(_03196_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07077_ (.I(_03196_),
    .Z(_03197_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07078_ (.A1(\u_cpu.rf_ram.memory[56][0] ),
    .A2(_03197_),
    .ZN(_03198_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07079_ (.A1(_03098_),
    .A2(_03197_),
    .B(_03198_),
    .ZN(_00461_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07080_ (.A1(\u_cpu.rf_ram.memory[56][1] ),
    .A2(_03197_),
    .ZN(_03199_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07081_ (.A1(_03102_),
    .A2(_03197_),
    .B(_03199_),
    .ZN(_00462_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07082_ (.A1(\u_cpu.rf_ram.memory[56][2] ),
    .A2(_03197_),
    .ZN(_03200_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07083_ (.A1(_03104_),
    .A2(_03197_),
    .B(_03200_),
    .ZN(_00463_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07084_ (.A1(\u_cpu.rf_ram.memory[56][3] ),
    .A2(_03197_),
    .ZN(_03201_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07085_ (.A1(_03106_),
    .A2(_03197_),
    .B(_03201_),
    .ZN(_00464_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07086_ (.A1(\u_cpu.rf_ram.memory[56][4] ),
    .A2(_03197_),
    .ZN(_03202_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07087_ (.A1(_03108_),
    .A2(_03197_),
    .B(_03202_),
    .ZN(_00465_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07088_ (.A1(\u_cpu.rf_ram.memory[56][5] ),
    .A2(_03197_),
    .ZN(_03203_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07089_ (.A1(_03110_),
    .A2(_03197_),
    .B(_03203_),
    .ZN(_00466_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07090_ (.A1(\u_cpu.rf_ram.memory[56][6] ),
    .A2(_03197_),
    .ZN(_03204_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07091_ (.A1(_03112_),
    .A2(_03197_),
    .B(_03204_),
    .ZN(_00467_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07092_ (.A1(\u_cpu.rf_ram.memory[56][7] ),
    .A2(_03197_),
    .ZN(_03205_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07093_ (.A1(_03114_),
    .A2(_03197_),
    .B(_03205_),
    .ZN(_00468_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07094_ (.A1(_02743_),
    .A2(_02827_),
    .ZN(_03206_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07095_ (.I(_03206_),
    .Z(_03207_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07096_ (.A1(\u_cpu.rf_ram.memory[55][0] ),
    .A2(_03207_),
    .ZN(_03208_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07097_ (.A1(_03098_),
    .A2(_03207_),
    .B(_03208_),
    .ZN(_00469_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07098_ (.A1(\u_cpu.rf_ram.memory[55][1] ),
    .A2(_03207_),
    .ZN(_03209_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07099_ (.A1(_03102_),
    .A2(_03207_),
    .B(_03209_),
    .ZN(_00470_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07100_ (.A1(\u_cpu.rf_ram.memory[55][2] ),
    .A2(_03207_),
    .ZN(_03210_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07101_ (.A1(_03104_),
    .A2(_03207_),
    .B(_03210_),
    .ZN(_00471_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07102_ (.A1(\u_cpu.rf_ram.memory[55][3] ),
    .A2(_03207_),
    .ZN(_03211_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07103_ (.A1(_03106_),
    .A2(_03207_),
    .B(_03211_),
    .ZN(_00472_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07104_ (.A1(\u_cpu.rf_ram.memory[55][4] ),
    .A2(_03207_),
    .ZN(_03212_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07105_ (.A1(_03108_),
    .A2(_03207_),
    .B(_03212_),
    .ZN(_00473_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07106_ (.A1(\u_cpu.rf_ram.memory[55][5] ),
    .A2(_03207_),
    .ZN(_03213_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07107_ (.A1(_03110_),
    .A2(_03207_),
    .B(_03213_),
    .ZN(_00474_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07108_ (.A1(\u_cpu.rf_ram.memory[55][6] ),
    .A2(_03207_),
    .ZN(_03214_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07109_ (.A1(_03112_),
    .A2(_03207_),
    .B(_03214_),
    .ZN(_00475_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07110_ (.A1(\u_cpu.rf_ram.memory[55][7] ),
    .A2(_03207_),
    .ZN(_03215_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07111_ (.A1(_03114_),
    .A2(_03207_),
    .B(_03215_),
    .ZN(_00476_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07112_ (.A1(_02827_),
    .A2(_03037_),
    .ZN(_03216_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07113_ (.I(_03216_),
    .Z(_03217_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07114_ (.A1(\u_cpu.rf_ram.memory[54][0] ),
    .A2(_03217_),
    .ZN(_03218_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07115_ (.A1(_03098_),
    .A2(_03217_),
    .B(_03218_),
    .ZN(_00477_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07116_ (.A1(\u_cpu.rf_ram.memory[54][1] ),
    .A2(_03217_),
    .ZN(_03219_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07117_ (.A1(_03102_),
    .A2(_03217_),
    .B(_03219_),
    .ZN(_00478_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07118_ (.A1(\u_cpu.rf_ram.memory[54][2] ),
    .A2(_03217_),
    .ZN(_03220_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07119_ (.A1(_03104_),
    .A2(_03217_),
    .B(_03220_),
    .ZN(_00479_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07120_ (.A1(\u_cpu.rf_ram.memory[54][3] ),
    .A2(_03217_),
    .ZN(_03221_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07121_ (.A1(_03106_),
    .A2(_03217_),
    .B(_03221_),
    .ZN(_00480_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07122_ (.A1(\u_cpu.rf_ram.memory[54][4] ),
    .A2(_03217_),
    .ZN(_03222_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07123_ (.A1(_03108_),
    .A2(_03217_),
    .B(_03222_),
    .ZN(_00481_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07124_ (.A1(\u_cpu.rf_ram.memory[54][5] ),
    .A2(_03217_),
    .ZN(_03223_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07125_ (.A1(_03110_),
    .A2(_03217_),
    .B(_03223_),
    .ZN(_00482_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07126_ (.A1(\u_cpu.rf_ram.memory[54][6] ),
    .A2(_03217_),
    .ZN(_03224_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07127_ (.A1(_03112_),
    .A2(_03217_),
    .B(_03224_),
    .ZN(_00483_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07128_ (.A1(\u_cpu.rf_ram.memory[54][7] ),
    .A2(_03217_),
    .ZN(_03225_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07129_ (.A1(_03114_),
    .A2(_03217_),
    .B(_03225_),
    .ZN(_00484_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07130_ (.A1(_02675_),
    .A2(_02827_),
    .ZN(_03226_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07131_ (.I(_03226_),
    .Z(_03227_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07132_ (.A1(\u_cpu.rf_ram.memory[53][0] ),
    .A2(_03227_),
    .ZN(_03228_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07133_ (.A1(_03098_),
    .A2(_03227_),
    .B(_03228_),
    .ZN(_00485_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07134_ (.A1(\u_cpu.rf_ram.memory[53][1] ),
    .A2(_03227_),
    .ZN(_03229_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07135_ (.A1(_03102_),
    .A2(_03227_),
    .B(_03229_),
    .ZN(_00486_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07136_ (.A1(\u_cpu.rf_ram.memory[53][2] ),
    .A2(_03227_),
    .ZN(_03230_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07137_ (.A1(_03104_),
    .A2(_03227_),
    .B(_03230_),
    .ZN(_00487_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07138_ (.A1(\u_cpu.rf_ram.memory[53][3] ),
    .A2(_03227_),
    .ZN(_03231_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07139_ (.A1(_03106_),
    .A2(_03227_),
    .B(_03231_),
    .ZN(_00488_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07140_ (.A1(\u_cpu.rf_ram.memory[53][4] ),
    .A2(_03227_),
    .ZN(_03232_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07141_ (.A1(_03108_),
    .A2(_03227_),
    .B(_03232_),
    .ZN(_00489_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07142_ (.A1(\u_cpu.rf_ram.memory[53][5] ),
    .A2(_03227_),
    .ZN(_03233_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07143_ (.A1(_03110_),
    .A2(_03227_),
    .B(_03233_),
    .ZN(_00490_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07144_ (.A1(\u_cpu.rf_ram.memory[53][6] ),
    .A2(_03227_),
    .ZN(_03234_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07145_ (.A1(_03112_),
    .A2(_03227_),
    .B(_03234_),
    .ZN(_00491_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07146_ (.A1(\u_cpu.rf_ram.memory[53][7] ),
    .A2(_03227_),
    .ZN(_03235_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07147_ (.A1(_03114_),
    .A2(_03227_),
    .B(_03235_),
    .ZN(_00492_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07148_ (.A1(_02717_),
    .A2(_02827_),
    .ZN(_03236_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07149_ (.I(_03236_),
    .Z(_03237_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07150_ (.A1(\u_cpu.rf_ram.memory[52][0] ),
    .A2(_03237_),
    .ZN(_03238_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07151_ (.A1(_03098_),
    .A2(_03237_),
    .B(_03238_),
    .ZN(_00493_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07152_ (.A1(\u_cpu.rf_ram.memory[52][1] ),
    .A2(_03237_),
    .ZN(_03239_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07153_ (.A1(_03102_),
    .A2(_03237_),
    .B(_03239_),
    .ZN(_00494_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07154_ (.A1(\u_cpu.rf_ram.memory[52][2] ),
    .A2(_03237_),
    .ZN(_03240_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07155_ (.A1(_03104_),
    .A2(_03237_),
    .B(_03240_),
    .ZN(_00495_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07156_ (.A1(\u_cpu.rf_ram.memory[52][3] ),
    .A2(_03237_),
    .ZN(_03241_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07157_ (.A1(_03106_),
    .A2(_03237_),
    .B(_03241_),
    .ZN(_00496_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07158_ (.A1(\u_cpu.rf_ram.memory[52][4] ),
    .A2(_03237_),
    .ZN(_03242_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07159_ (.A1(_03108_),
    .A2(_03237_),
    .B(_03242_),
    .ZN(_00497_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07160_ (.A1(\u_cpu.rf_ram.memory[52][5] ),
    .A2(_03237_),
    .ZN(_03243_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07161_ (.A1(_03110_),
    .A2(_03237_),
    .B(_03243_),
    .ZN(_00498_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07162_ (.A1(\u_cpu.rf_ram.memory[52][6] ),
    .A2(_03237_),
    .ZN(_03244_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07163_ (.A1(_03112_),
    .A2(_03237_),
    .B(_03244_),
    .ZN(_00499_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07164_ (.A1(\u_cpu.rf_ram.memory[52][7] ),
    .A2(_03237_),
    .ZN(_03245_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07165_ (.A1(_03114_),
    .A2(_03237_),
    .B(_03245_),
    .ZN(_00500_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _07166_ (.A1(_02731_),
    .A2(_02838_),
    .Z(_03246_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07167_ (.I(_03246_),
    .Z(_03247_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07168_ (.A1(\u_cpu.rf_ram.memory[9][0] ),
    .A2(_03247_),
    .ZN(_03248_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07169_ (.A1(_02632_),
    .A2(_03247_),
    .B(_03248_),
    .ZN(_00501_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07170_ (.A1(\u_cpu.rf_ram.memory[9][1] ),
    .A2(_03247_),
    .ZN(_03249_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07171_ (.A1(_02637_),
    .A2(_03247_),
    .B(_03249_),
    .ZN(_00502_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07172_ (.A1(\u_cpu.rf_ram.memory[9][2] ),
    .A2(_03247_),
    .ZN(_03250_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07173_ (.A1(_02642_),
    .A2(_03247_),
    .B(_03250_),
    .ZN(_00503_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07174_ (.A1(\u_cpu.rf_ram.memory[9][3] ),
    .A2(_03247_),
    .ZN(_03251_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07175_ (.A1(_02647_),
    .A2(_03247_),
    .B(_03251_),
    .ZN(_00504_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07176_ (.A1(\u_cpu.rf_ram.memory[9][4] ),
    .A2(_03247_),
    .ZN(_03252_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07177_ (.A1(_02652_),
    .A2(_03247_),
    .B(_03252_),
    .ZN(_00505_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07178_ (.A1(\u_cpu.rf_ram.memory[9][5] ),
    .A2(_03247_),
    .ZN(_03253_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07179_ (.A1(_02657_),
    .A2(_03247_),
    .B(_03253_),
    .ZN(_00506_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07180_ (.A1(\u_cpu.rf_ram.memory[9][6] ),
    .A2(_03247_),
    .ZN(_03254_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07181_ (.A1(_02662_),
    .A2(_03247_),
    .B(_03254_),
    .ZN(_00507_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07182_ (.A1(\u_cpu.rf_ram.memory[9][7] ),
    .A2(_03247_),
    .ZN(_03255_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07183_ (.A1(_02667_),
    .A2(_03247_),
    .B(_03255_),
    .ZN(_00508_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07184_ (.A1(_02731_),
    .A2(_02870_),
    .ZN(_03256_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07185_ (.I(_03256_),
    .ZN(_03257_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07186_ (.A1(\u_cpu.rf_ram.memory[15][0] ),
    .A2(_03257_),
    .ZN(_03258_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07187_ (.A1(_02632_),
    .A2(_03257_),
    .B(_03258_),
    .ZN(_00509_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07188_ (.A1(\u_cpu.rf_ram.memory[15][1] ),
    .A2(_03257_),
    .ZN(_03259_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07189_ (.A1(_02637_),
    .A2(_03257_),
    .B(_03259_),
    .ZN(_00510_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07190_ (.A1(\u_cpu.rf_ram.memory[15][2] ),
    .A2(_03257_),
    .ZN(_03260_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07191_ (.A1(_02642_),
    .A2(_03257_),
    .B(_03260_),
    .ZN(_00511_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07192_ (.A1(\u_cpu.rf_ram.memory[15][3] ),
    .A2(_03257_),
    .ZN(_03261_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07193_ (.A1(_02647_),
    .A2(_03257_),
    .B(_03261_),
    .ZN(_00512_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07194_ (.A1(\u_cpu.rf_ram.memory[15][4] ),
    .A2(_03257_),
    .ZN(_03262_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07195_ (.A1(_02652_),
    .A2(_03257_),
    .B(_03262_),
    .ZN(_00513_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07196_ (.A1(\u_cpu.rf_ram.memory[15][5] ),
    .A2(_03257_),
    .ZN(_03263_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07197_ (.A1(_02657_),
    .A2(_03257_),
    .B(_03263_),
    .ZN(_00514_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07198_ (.A1(\u_cpu.rf_ram.memory[15][6] ),
    .A2(_03257_),
    .ZN(_03264_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07199_ (.A1(_02662_),
    .A2(_03257_),
    .B(_03264_),
    .ZN(_00515_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07200_ (.A1(\u_cpu.rf_ram.memory[15][7] ),
    .A2(_03257_),
    .ZN(_03265_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07201_ (.A1(_02667_),
    .A2(_03257_),
    .B(_03265_),
    .ZN(_00516_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07202_ (.A1(_02766_),
    .A2(_02976_),
    .ZN(_03266_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07203_ (.I(_03266_),
    .Z(_03267_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07204_ (.A1(\u_cpu.rf_ram.memory[142][0] ),
    .A2(_03267_),
    .ZN(_03268_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07205_ (.A1(_03098_),
    .A2(_03267_),
    .B(_03268_),
    .ZN(_00517_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07206_ (.A1(\u_cpu.rf_ram.memory[142][1] ),
    .A2(_03267_),
    .ZN(_03269_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07207_ (.A1(_03102_),
    .A2(_03267_),
    .B(_03269_),
    .ZN(_00518_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07208_ (.A1(\u_cpu.rf_ram.memory[142][2] ),
    .A2(_03267_),
    .ZN(_03270_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07209_ (.A1(_03104_),
    .A2(_03267_),
    .B(_03270_),
    .ZN(_00519_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07210_ (.A1(\u_cpu.rf_ram.memory[142][3] ),
    .A2(_03267_),
    .ZN(_03271_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07211_ (.A1(_03106_),
    .A2(_03267_),
    .B(_03271_),
    .ZN(_00520_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07212_ (.A1(\u_cpu.rf_ram.memory[142][4] ),
    .A2(_03267_),
    .ZN(_03272_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07213_ (.A1(_03108_),
    .A2(_03267_),
    .B(_03272_),
    .ZN(_00521_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07214_ (.A1(\u_cpu.rf_ram.memory[142][5] ),
    .A2(_03267_),
    .ZN(_03273_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07215_ (.A1(_03110_),
    .A2(_03267_),
    .B(_03273_),
    .ZN(_00522_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07216_ (.A1(\u_cpu.rf_ram.memory[142][6] ),
    .A2(_03267_),
    .ZN(_03274_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07217_ (.A1(_03112_),
    .A2(_03267_),
    .B(_03274_),
    .ZN(_00523_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07218_ (.A1(\u_cpu.rf_ram.memory[142][7] ),
    .A2(_03267_),
    .ZN(_03275_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07219_ (.A1(_03114_),
    .A2(_03267_),
    .B(_03275_),
    .ZN(_00524_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07220_ (.A1(_02803_),
    .A2(_02976_),
    .ZN(_03276_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07221_ (.I(_03276_),
    .Z(_03277_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07222_ (.A1(\u_cpu.rf_ram.memory[141][0] ),
    .A2(_03277_),
    .ZN(_03278_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07223_ (.A1(_03098_),
    .A2(_03277_),
    .B(_03278_),
    .ZN(_00525_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07224_ (.A1(\u_cpu.rf_ram.memory[141][1] ),
    .A2(_03277_),
    .ZN(_03279_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07225_ (.A1(_03102_),
    .A2(_03277_),
    .B(_03279_),
    .ZN(_00526_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07226_ (.A1(\u_cpu.rf_ram.memory[141][2] ),
    .A2(_03277_),
    .ZN(_03280_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07227_ (.A1(_03104_),
    .A2(_03277_),
    .B(_03280_),
    .ZN(_00527_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07228_ (.A1(\u_cpu.rf_ram.memory[141][3] ),
    .A2(_03277_),
    .ZN(_03281_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07229_ (.A1(_03106_),
    .A2(_03277_),
    .B(_03281_),
    .ZN(_00528_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07230_ (.A1(\u_cpu.rf_ram.memory[141][4] ),
    .A2(_03277_),
    .ZN(_03282_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07231_ (.A1(_03108_),
    .A2(_03277_),
    .B(_03282_),
    .ZN(_00529_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07232_ (.A1(\u_cpu.rf_ram.memory[141][5] ),
    .A2(_03277_),
    .ZN(_03283_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07233_ (.A1(_03110_),
    .A2(_03277_),
    .B(_03283_),
    .ZN(_00530_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07234_ (.A1(\u_cpu.rf_ram.memory[141][6] ),
    .A2(_03277_),
    .ZN(_03284_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07235_ (.A1(_03112_),
    .A2(_03277_),
    .B(_03284_),
    .ZN(_00531_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07236_ (.A1(\u_cpu.rf_ram.memory[141][7] ),
    .A2(_03277_),
    .ZN(_03285_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07237_ (.A1(_03114_),
    .A2(_03277_),
    .B(_03285_),
    .ZN(_00532_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07238_ (.A1(_02814_),
    .A2(_02976_),
    .ZN(_03286_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07239_ (.I(_03286_),
    .Z(_03287_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07240_ (.A1(\u_cpu.rf_ram.memory[140][0] ),
    .A2(_03287_),
    .ZN(_03288_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07241_ (.A1(_03098_),
    .A2(_03287_),
    .B(_03288_),
    .ZN(_00533_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07242_ (.A1(\u_cpu.rf_ram.memory[140][1] ),
    .A2(_03287_),
    .ZN(_03289_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07243_ (.A1(_03102_),
    .A2(_03287_),
    .B(_03289_),
    .ZN(_00534_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07244_ (.A1(\u_cpu.rf_ram.memory[140][2] ),
    .A2(_03287_),
    .ZN(_03290_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07245_ (.A1(_03104_),
    .A2(_03287_),
    .B(_03290_),
    .ZN(_00535_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07246_ (.A1(\u_cpu.rf_ram.memory[140][3] ),
    .A2(_03287_),
    .ZN(_03291_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07247_ (.A1(_03106_),
    .A2(_03287_),
    .B(_03291_),
    .ZN(_00536_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07248_ (.A1(\u_cpu.rf_ram.memory[140][4] ),
    .A2(_03287_),
    .ZN(_03292_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07249_ (.A1(_03108_),
    .A2(_03287_),
    .B(_03292_),
    .ZN(_00537_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07250_ (.A1(\u_cpu.rf_ram.memory[140][5] ),
    .A2(_03287_),
    .ZN(_03293_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07251_ (.A1(_03110_),
    .A2(_03287_),
    .B(_03293_),
    .ZN(_00538_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07252_ (.A1(\u_cpu.rf_ram.memory[140][6] ),
    .A2(_03287_),
    .ZN(_03294_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07253_ (.A1(_03112_),
    .A2(_03287_),
    .B(_03294_),
    .ZN(_00539_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07254_ (.A1(\u_cpu.rf_ram.memory[140][7] ),
    .A2(_03287_),
    .ZN(_03295_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07255_ (.A1(_03114_),
    .A2(_03287_),
    .B(_03295_),
    .ZN(_00540_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07256_ (.A1(_02731_),
    .A2(_02803_),
    .ZN(_03296_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07257_ (.I(_03296_),
    .ZN(_03297_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07258_ (.A1(\u_cpu.rf_ram.memory[13][0] ),
    .A2(_03297_),
    .ZN(_03298_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07259_ (.A1(_02632_),
    .A2(_03297_),
    .B(_03298_),
    .ZN(_00541_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07260_ (.A1(\u_cpu.rf_ram.memory[13][1] ),
    .A2(_03297_),
    .ZN(_03299_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07261_ (.A1(_02637_),
    .A2(_03297_),
    .B(_03299_),
    .ZN(_00542_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07262_ (.A1(\u_cpu.rf_ram.memory[13][2] ),
    .A2(_03297_),
    .ZN(_03300_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07263_ (.A1(_02642_),
    .A2(_03297_),
    .B(_03300_),
    .ZN(_00543_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07264_ (.A1(\u_cpu.rf_ram.memory[13][3] ),
    .A2(_03297_),
    .ZN(_03301_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07265_ (.A1(_02647_),
    .A2(_03297_),
    .B(_03301_),
    .ZN(_00544_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07266_ (.A1(\u_cpu.rf_ram.memory[13][4] ),
    .A2(_03297_),
    .ZN(_03302_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07267_ (.A1(_02652_),
    .A2(_03297_),
    .B(_03302_),
    .ZN(_00545_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07268_ (.A1(\u_cpu.rf_ram.memory[13][5] ),
    .A2(_03297_),
    .ZN(_03303_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07269_ (.A1(_02657_),
    .A2(_03297_),
    .B(_03303_),
    .ZN(_00546_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07270_ (.A1(\u_cpu.rf_ram.memory[13][6] ),
    .A2(_03297_),
    .ZN(_03304_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07271_ (.A1(_02662_),
    .A2(_03297_),
    .B(_03304_),
    .ZN(_00547_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07272_ (.A1(\u_cpu.rf_ram.memory[13][7] ),
    .A2(_03297_),
    .ZN(_03305_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07273_ (.A1(_02667_),
    .A2(_03297_),
    .B(_03305_),
    .ZN(_00548_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07274_ (.I(_02631_),
    .Z(_03306_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07275_ (.A1(_02768_),
    .A2(_02954_),
    .ZN(_03307_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07276_ (.I(_03307_),
    .Z(_03308_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07277_ (.A1(\u_cpu.rf_ram.memory[72][0] ),
    .A2(_03308_),
    .ZN(_03309_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07278_ (.A1(_03306_),
    .A2(_03308_),
    .B(_03309_),
    .ZN(_00549_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07279_ (.I(_02636_),
    .Z(_03310_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07280_ (.A1(\u_cpu.rf_ram.memory[72][1] ),
    .A2(_03308_),
    .ZN(_03311_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07281_ (.A1(_03310_),
    .A2(_03308_),
    .B(_03311_),
    .ZN(_00550_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07282_ (.I(_02641_),
    .Z(_03312_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07283_ (.A1(\u_cpu.rf_ram.memory[72][2] ),
    .A2(_03308_),
    .ZN(_03313_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07284_ (.A1(_03312_),
    .A2(_03308_),
    .B(_03313_),
    .ZN(_00551_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07285_ (.I(_02646_),
    .Z(_03314_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07286_ (.A1(\u_cpu.rf_ram.memory[72][3] ),
    .A2(_03308_),
    .ZN(_03315_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07287_ (.A1(_03314_),
    .A2(_03308_),
    .B(_03315_),
    .ZN(_00552_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07288_ (.I(_02651_),
    .Z(_03316_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07289_ (.A1(\u_cpu.rf_ram.memory[72][4] ),
    .A2(_03308_),
    .ZN(_03317_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07290_ (.A1(_03316_),
    .A2(_03308_),
    .B(_03317_),
    .ZN(_00553_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07291_ (.I(_02656_),
    .Z(_03318_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07292_ (.A1(\u_cpu.rf_ram.memory[72][5] ),
    .A2(_03308_),
    .ZN(_03319_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07293_ (.A1(_03318_),
    .A2(_03308_),
    .B(_03319_),
    .ZN(_00554_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07294_ (.I(_02661_),
    .Z(_03320_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07295_ (.A1(\u_cpu.rf_ram.memory[72][6] ),
    .A2(_03308_),
    .ZN(_03321_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07296_ (.A1(_03320_),
    .A2(_03308_),
    .B(_03321_),
    .ZN(_00555_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07297_ (.I(_02666_),
    .Z(_03322_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07298_ (.A1(\u_cpu.rf_ram.memory[72][7] ),
    .A2(_03308_),
    .ZN(_03323_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07299_ (.A1(_03322_),
    .A2(_03308_),
    .B(_03323_),
    .ZN(_00556_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07300_ (.A1(_02768_),
    .A2(_02838_),
    .ZN(_03324_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07301_ (.I(_03324_),
    .Z(_03325_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07302_ (.A1(\u_cpu.rf_ram.memory[73][0] ),
    .A2(_03325_),
    .ZN(_03326_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07303_ (.A1(_03306_),
    .A2(_03325_),
    .B(_03326_),
    .ZN(_00557_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07304_ (.A1(\u_cpu.rf_ram.memory[73][1] ),
    .A2(_03325_),
    .ZN(_03327_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07305_ (.A1(_03310_),
    .A2(_03325_),
    .B(_03327_),
    .ZN(_00558_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07306_ (.A1(\u_cpu.rf_ram.memory[73][2] ),
    .A2(_03325_),
    .ZN(_03328_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07307_ (.A1(_03312_),
    .A2(_03325_),
    .B(_03328_),
    .ZN(_00559_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07308_ (.A1(\u_cpu.rf_ram.memory[73][3] ),
    .A2(_03325_),
    .ZN(_03329_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07309_ (.A1(_03314_),
    .A2(_03325_),
    .B(_03329_),
    .ZN(_00560_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07310_ (.A1(\u_cpu.rf_ram.memory[73][4] ),
    .A2(_03325_),
    .ZN(_03330_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07311_ (.A1(_03316_),
    .A2(_03325_),
    .B(_03330_),
    .ZN(_00561_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07312_ (.A1(\u_cpu.rf_ram.memory[73][5] ),
    .A2(_03325_),
    .ZN(_03331_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07313_ (.A1(_03318_),
    .A2(_03325_),
    .B(_03331_),
    .ZN(_00562_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07314_ (.A1(\u_cpu.rf_ram.memory[73][6] ),
    .A2(_03325_),
    .ZN(_03332_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07315_ (.A1(_03320_),
    .A2(_03325_),
    .B(_03332_),
    .ZN(_00563_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07316_ (.A1(\u_cpu.rf_ram.memory[73][7] ),
    .A2(_03325_),
    .ZN(_03333_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07317_ (.A1(_03322_),
    .A2(_03325_),
    .B(_03333_),
    .ZN(_00564_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07318_ (.A1(_02743_),
    .A2(_02768_),
    .ZN(_03334_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07319_ (.I(_03334_),
    .Z(_03335_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07320_ (.A1(\u_cpu.rf_ram.memory[71][0] ),
    .A2(_03335_),
    .ZN(_03336_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07321_ (.A1(_03306_),
    .A2(_03335_),
    .B(_03336_),
    .ZN(_00565_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07322_ (.A1(\u_cpu.rf_ram.memory[71][1] ),
    .A2(_03335_),
    .ZN(_03337_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07323_ (.A1(_03310_),
    .A2(_03335_),
    .B(_03337_),
    .ZN(_00566_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07324_ (.A1(\u_cpu.rf_ram.memory[71][2] ),
    .A2(_03335_),
    .ZN(_03338_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07325_ (.A1(_03312_),
    .A2(_03335_),
    .B(_03338_),
    .ZN(_00567_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07326_ (.A1(\u_cpu.rf_ram.memory[71][3] ),
    .A2(_03335_),
    .ZN(_03339_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07327_ (.A1(_03314_),
    .A2(_03335_),
    .B(_03339_),
    .ZN(_00568_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07328_ (.A1(\u_cpu.rf_ram.memory[71][4] ),
    .A2(_03335_),
    .ZN(_03340_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07329_ (.A1(_03316_),
    .A2(_03335_),
    .B(_03340_),
    .ZN(_00569_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07330_ (.A1(\u_cpu.rf_ram.memory[71][5] ),
    .A2(_03335_),
    .ZN(_03341_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07331_ (.A1(_03318_),
    .A2(_03335_),
    .B(_03341_),
    .ZN(_00570_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07332_ (.A1(\u_cpu.rf_ram.memory[71][6] ),
    .A2(_03335_),
    .ZN(_03342_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07333_ (.A1(_03320_),
    .A2(_03335_),
    .B(_03342_),
    .ZN(_00571_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07334_ (.A1(\u_cpu.rf_ram.memory[71][7] ),
    .A2(_03335_),
    .ZN(_03343_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07335_ (.A1(_03322_),
    .A2(_03335_),
    .B(_03343_),
    .ZN(_00572_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07336_ (.A1(_02768_),
    .A2(_03037_),
    .ZN(_03344_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07337_ (.I(_03344_),
    .Z(_03345_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07338_ (.A1(\u_cpu.rf_ram.memory[70][0] ),
    .A2(_03345_),
    .ZN(_03346_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07339_ (.A1(_03306_),
    .A2(_03345_),
    .B(_03346_),
    .ZN(_00573_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07340_ (.A1(\u_cpu.rf_ram.memory[70][1] ),
    .A2(_03345_),
    .ZN(_03347_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07341_ (.A1(_03310_),
    .A2(_03345_),
    .B(_03347_),
    .ZN(_00574_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07342_ (.A1(\u_cpu.rf_ram.memory[70][2] ),
    .A2(_03345_),
    .ZN(_03348_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07343_ (.A1(_03312_),
    .A2(_03345_),
    .B(_03348_),
    .ZN(_00575_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07344_ (.A1(\u_cpu.rf_ram.memory[70][3] ),
    .A2(_03345_),
    .ZN(_03349_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07345_ (.A1(_03314_),
    .A2(_03345_),
    .B(_03349_),
    .ZN(_00576_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07346_ (.A1(\u_cpu.rf_ram.memory[70][4] ),
    .A2(_03345_),
    .ZN(_03350_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07347_ (.A1(_03316_),
    .A2(_03345_),
    .B(_03350_),
    .ZN(_00577_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07348_ (.A1(\u_cpu.rf_ram.memory[70][5] ),
    .A2(_03345_),
    .ZN(_03351_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07349_ (.A1(_03318_),
    .A2(_03345_),
    .B(_03351_),
    .ZN(_00578_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07350_ (.A1(\u_cpu.rf_ram.memory[70][6] ),
    .A2(_03345_),
    .ZN(_03352_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07351_ (.A1(_03320_),
    .A2(_03345_),
    .B(_03352_),
    .ZN(_00579_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07352_ (.A1(\u_cpu.rf_ram.memory[70][7] ),
    .A2(_03345_),
    .ZN(_03353_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07353_ (.A1(_03322_),
    .A2(_03345_),
    .B(_03353_),
    .ZN(_00580_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07354_ (.A1(_02870_),
    .A2(_02976_),
    .ZN(_03354_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07355_ (.I(_03354_),
    .Z(_03355_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07356_ (.A1(\u_cpu.rf_ram.memory[143][0] ),
    .A2(_03355_),
    .ZN(_03356_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07357_ (.A1(_03306_),
    .A2(_03355_),
    .B(_03356_),
    .ZN(_00581_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07358_ (.A1(\u_cpu.rf_ram.memory[143][1] ),
    .A2(_03355_),
    .ZN(_03357_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07359_ (.A1(_03310_),
    .A2(_03355_),
    .B(_03357_),
    .ZN(_00582_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07360_ (.A1(\u_cpu.rf_ram.memory[143][2] ),
    .A2(_03355_),
    .ZN(_03358_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07361_ (.A1(_03312_),
    .A2(_03355_),
    .B(_03358_),
    .ZN(_00583_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07362_ (.A1(\u_cpu.rf_ram.memory[143][3] ),
    .A2(_03355_),
    .ZN(_03359_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07363_ (.A1(_03314_),
    .A2(_03355_),
    .B(_03359_),
    .ZN(_00584_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07364_ (.A1(\u_cpu.rf_ram.memory[143][4] ),
    .A2(_03355_),
    .ZN(_03360_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07365_ (.A1(_03316_),
    .A2(_03355_),
    .B(_03360_),
    .ZN(_00585_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07366_ (.A1(\u_cpu.rf_ram.memory[143][5] ),
    .A2(_03355_),
    .ZN(_03361_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07367_ (.A1(_03318_),
    .A2(_03355_),
    .B(_03361_),
    .ZN(_00586_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07368_ (.A1(\u_cpu.rf_ram.memory[143][6] ),
    .A2(_03355_),
    .ZN(_03362_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07369_ (.A1(_03320_),
    .A2(_03355_),
    .B(_03362_),
    .ZN(_00587_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07370_ (.A1(\u_cpu.rf_ram.memory[143][7] ),
    .A2(_03355_),
    .ZN(_03363_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07371_ (.A1(_03322_),
    .A2(_03355_),
    .B(_03363_),
    .ZN(_00588_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07372_ (.A1(_02731_),
    .A2(_02766_),
    .ZN(_03364_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07373_ (.I(_03364_),
    .ZN(_03365_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07374_ (.A1(\u_cpu.rf_ram.memory[14][0] ),
    .A2(_03365_),
    .ZN(_03366_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07375_ (.A1(_02632_),
    .A2(_03365_),
    .B(_03366_),
    .ZN(_00589_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07376_ (.A1(\u_cpu.rf_ram.memory[14][1] ),
    .A2(_03365_),
    .ZN(_03367_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07377_ (.A1(_02637_),
    .A2(_03365_),
    .B(_03367_),
    .ZN(_00590_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07378_ (.A1(\u_cpu.rf_ram.memory[14][2] ),
    .A2(_03365_),
    .ZN(_03368_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07379_ (.A1(_02642_),
    .A2(_03365_),
    .B(_03368_),
    .ZN(_00591_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07380_ (.A1(\u_cpu.rf_ram.memory[14][3] ),
    .A2(_03365_),
    .ZN(_03369_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07381_ (.A1(_02647_),
    .A2(_03365_),
    .B(_03369_),
    .ZN(_00592_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07382_ (.A1(\u_cpu.rf_ram.memory[14][4] ),
    .A2(_03365_),
    .ZN(_03370_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07383_ (.A1(_02652_),
    .A2(_03365_),
    .B(_03370_),
    .ZN(_00593_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07384_ (.A1(\u_cpu.rf_ram.memory[14][5] ),
    .A2(_03365_),
    .ZN(_03371_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07385_ (.A1(_02657_),
    .A2(_03365_),
    .B(_03371_),
    .ZN(_00594_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07386_ (.A1(\u_cpu.rf_ram.memory[14][6] ),
    .A2(_03365_),
    .ZN(_03372_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07387_ (.A1(_02662_),
    .A2(_03365_),
    .B(_03372_),
    .ZN(_00595_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07388_ (.A1(\u_cpu.rf_ram.memory[14][7] ),
    .A2(_03365_),
    .ZN(_03373_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07389_ (.A1(_02667_),
    .A2(_03365_),
    .B(_03373_),
    .ZN(_00596_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07390_ (.A1(_02780_),
    .A2(_02976_),
    .ZN(_03374_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07391_ (.I(_03374_),
    .Z(_03375_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07392_ (.A1(\u_cpu.rf_ram.memory[138][0] ),
    .A2(_03375_),
    .ZN(_03376_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07393_ (.A1(_03306_),
    .A2(_03375_),
    .B(_03376_),
    .ZN(_00597_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07394_ (.A1(\u_cpu.rf_ram.memory[138][1] ),
    .A2(_03375_),
    .ZN(_03377_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07395_ (.A1(_03310_),
    .A2(_03375_),
    .B(_03377_),
    .ZN(_00598_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07396_ (.A1(\u_cpu.rf_ram.memory[138][2] ),
    .A2(_03375_),
    .ZN(_03378_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07397_ (.A1(_03312_),
    .A2(_03375_),
    .B(_03378_),
    .ZN(_00599_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07398_ (.A1(\u_cpu.rf_ram.memory[138][3] ),
    .A2(_03375_),
    .ZN(_03379_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07399_ (.A1(_03314_),
    .A2(_03375_),
    .B(_03379_),
    .ZN(_00600_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07400_ (.A1(\u_cpu.rf_ram.memory[138][4] ),
    .A2(_03375_),
    .ZN(_03380_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07401_ (.A1(_03316_),
    .A2(_03375_),
    .B(_03380_),
    .ZN(_00601_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07402_ (.A1(\u_cpu.rf_ram.memory[138][5] ),
    .A2(_03375_),
    .ZN(_03381_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07403_ (.A1(_03318_),
    .A2(_03375_),
    .B(_03381_),
    .ZN(_00602_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07404_ (.A1(\u_cpu.rf_ram.memory[138][6] ),
    .A2(_03375_),
    .ZN(_03382_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07405_ (.A1(_03320_),
    .A2(_03375_),
    .B(_03382_),
    .ZN(_00603_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07406_ (.A1(\u_cpu.rf_ram.memory[138][7] ),
    .A2(_03375_),
    .ZN(_03383_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07407_ (.A1(_03322_),
    .A2(_03375_),
    .B(_03383_),
    .ZN(_00604_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07408_ (.A1(_02743_),
    .A2(_02782_),
    .ZN(_03384_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07409_ (.I(_03384_),
    .Z(_03385_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07410_ (.A1(\u_cpu.rf_ram.memory[39][0] ),
    .A2(_03385_),
    .ZN(_03386_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07411_ (.A1(_03306_),
    .A2(_03385_),
    .B(_03386_),
    .ZN(_00605_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07412_ (.A1(\u_cpu.rf_ram.memory[39][1] ),
    .A2(_03385_),
    .ZN(_03387_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07413_ (.A1(_03310_),
    .A2(_03385_),
    .B(_03387_),
    .ZN(_00606_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07414_ (.A1(\u_cpu.rf_ram.memory[39][2] ),
    .A2(_03385_),
    .ZN(_03388_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07415_ (.A1(_03312_),
    .A2(_03385_),
    .B(_03388_),
    .ZN(_00607_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07416_ (.A1(\u_cpu.rf_ram.memory[39][3] ),
    .A2(_03385_),
    .ZN(_03389_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07417_ (.A1(_03314_),
    .A2(_03385_),
    .B(_03389_),
    .ZN(_00608_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07418_ (.A1(\u_cpu.rf_ram.memory[39][4] ),
    .A2(_03385_),
    .ZN(_03390_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07419_ (.A1(_03316_),
    .A2(_03385_),
    .B(_03390_),
    .ZN(_00609_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07420_ (.A1(\u_cpu.rf_ram.memory[39][5] ),
    .A2(_03385_),
    .ZN(_03391_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07421_ (.A1(_03318_),
    .A2(_03385_),
    .B(_03391_),
    .ZN(_00610_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07422_ (.A1(\u_cpu.rf_ram.memory[39][6] ),
    .A2(_03385_),
    .ZN(_03392_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07423_ (.A1(_03320_),
    .A2(_03385_),
    .B(_03392_),
    .ZN(_00611_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07424_ (.A1(\u_cpu.rf_ram.memory[39][7] ),
    .A2(_03385_),
    .ZN(_03393_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07425_ (.A1(_03322_),
    .A2(_03385_),
    .B(_03393_),
    .ZN(_00612_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07426_ (.A1(_02838_),
    .A2(_02976_),
    .ZN(_03394_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07427_ (.I(_03394_),
    .Z(_03395_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07428_ (.A1(\u_cpu.rf_ram.memory[137][0] ),
    .A2(_03395_),
    .ZN(_03396_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07429_ (.A1(_03306_),
    .A2(_03395_),
    .B(_03396_),
    .ZN(_00613_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07430_ (.A1(\u_cpu.rf_ram.memory[137][1] ),
    .A2(_03395_),
    .ZN(_03397_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07431_ (.A1(_03310_),
    .A2(_03395_),
    .B(_03397_),
    .ZN(_00614_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07432_ (.A1(\u_cpu.rf_ram.memory[137][2] ),
    .A2(_03395_),
    .ZN(_03398_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07433_ (.A1(_03312_),
    .A2(_03395_),
    .B(_03398_),
    .ZN(_00615_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07434_ (.A1(\u_cpu.rf_ram.memory[137][3] ),
    .A2(_03395_),
    .ZN(_03399_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07435_ (.A1(_03314_),
    .A2(_03395_),
    .B(_03399_),
    .ZN(_00616_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07436_ (.A1(\u_cpu.rf_ram.memory[137][4] ),
    .A2(_03395_),
    .ZN(_03400_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07437_ (.A1(_03316_),
    .A2(_03395_),
    .B(_03400_),
    .ZN(_00617_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07438_ (.A1(\u_cpu.rf_ram.memory[137][5] ),
    .A2(_03395_),
    .ZN(_03401_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07439_ (.A1(_03318_),
    .A2(_03395_),
    .B(_03401_),
    .ZN(_00618_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07440_ (.A1(\u_cpu.rf_ram.memory[137][6] ),
    .A2(_03395_),
    .ZN(_03402_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07441_ (.A1(_03320_),
    .A2(_03395_),
    .B(_03402_),
    .ZN(_00619_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07442_ (.A1(\u_cpu.rf_ram.memory[137][7] ),
    .A2(_03395_),
    .ZN(_03403_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07443_ (.A1(_03322_),
    .A2(_03395_),
    .B(_03403_),
    .ZN(_00620_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07444_ (.A1(_02695_),
    .A2(_02827_),
    .ZN(_03404_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07445_ (.I(_03404_),
    .Z(_03405_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07446_ (.A1(\u_cpu.rf_ram.memory[49][0] ),
    .A2(_03405_),
    .ZN(_03406_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07447_ (.A1(_03306_),
    .A2(_03405_),
    .B(_03406_),
    .ZN(_00621_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07448_ (.A1(\u_cpu.rf_ram.memory[49][1] ),
    .A2(_03405_),
    .ZN(_03407_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07449_ (.A1(_03310_),
    .A2(_03405_),
    .B(_03407_),
    .ZN(_00622_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07450_ (.A1(\u_cpu.rf_ram.memory[49][2] ),
    .A2(_03405_),
    .ZN(_03408_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07451_ (.A1(_03312_),
    .A2(_03405_),
    .B(_03408_),
    .ZN(_00623_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07452_ (.A1(\u_cpu.rf_ram.memory[49][3] ),
    .A2(_03405_),
    .ZN(_03409_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07453_ (.A1(_03314_),
    .A2(_03405_),
    .B(_03409_),
    .ZN(_00624_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07454_ (.A1(\u_cpu.rf_ram.memory[49][4] ),
    .A2(_03405_),
    .ZN(_03410_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07455_ (.A1(_03316_),
    .A2(_03405_),
    .B(_03410_),
    .ZN(_00625_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07456_ (.A1(\u_cpu.rf_ram.memory[49][5] ),
    .A2(_03405_),
    .ZN(_03411_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07457_ (.A1(_03318_),
    .A2(_03405_),
    .B(_03411_),
    .ZN(_00626_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07458_ (.A1(\u_cpu.rf_ram.memory[49][6] ),
    .A2(_03405_),
    .ZN(_03412_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07459_ (.A1(_03320_),
    .A2(_03405_),
    .B(_03412_),
    .ZN(_00627_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07460_ (.A1(\u_cpu.rf_ram.memory[49][7] ),
    .A2(_03405_),
    .ZN(_03413_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07461_ (.A1(_03322_),
    .A2(_03405_),
    .B(_03413_),
    .ZN(_00628_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07462_ (.A1(_02954_),
    .A2(_02976_),
    .ZN(_03414_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07463_ (.I(_03414_),
    .Z(_03415_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07464_ (.A1(\u_cpu.rf_ram.memory[136][0] ),
    .A2(_03415_),
    .ZN(_03416_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07465_ (.A1(_03306_),
    .A2(_03415_),
    .B(_03416_),
    .ZN(_00629_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07466_ (.A1(\u_cpu.rf_ram.memory[136][1] ),
    .A2(_03415_),
    .ZN(_03417_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07467_ (.A1(_03310_),
    .A2(_03415_),
    .B(_03417_),
    .ZN(_00630_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07468_ (.A1(\u_cpu.rf_ram.memory[136][2] ),
    .A2(_03415_),
    .ZN(_03418_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07469_ (.A1(_03312_),
    .A2(_03415_),
    .B(_03418_),
    .ZN(_00631_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07470_ (.A1(\u_cpu.rf_ram.memory[136][3] ),
    .A2(_03415_),
    .ZN(_03419_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07471_ (.A1(_03314_),
    .A2(_03415_),
    .B(_03419_),
    .ZN(_00632_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07472_ (.A1(\u_cpu.rf_ram.memory[136][4] ),
    .A2(_03415_),
    .ZN(_03420_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07473_ (.A1(_03316_),
    .A2(_03415_),
    .B(_03420_),
    .ZN(_00633_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07474_ (.A1(\u_cpu.rf_ram.memory[136][5] ),
    .A2(_03415_),
    .ZN(_03421_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07475_ (.A1(_03318_),
    .A2(_03415_),
    .B(_03421_),
    .ZN(_00634_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07476_ (.A1(\u_cpu.rf_ram.memory[136][6] ),
    .A2(_03415_),
    .ZN(_03422_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07477_ (.A1(_03320_),
    .A2(_03415_),
    .B(_03422_),
    .ZN(_00635_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07478_ (.A1(\u_cpu.rf_ram.memory[136][7] ),
    .A2(_03415_),
    .ZN(_03423_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07479_ (.A1(_03322_),
    .A2(_03415_),
    .B(_03423_),
    .ZN(_00636_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07480_ (.A1(_02743_),
    .A2(_02976_),
    .ZN(_03424_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07481_ (.I(_03424_),
    .Z(_03425_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07482_ (.A1(\u_cpu.rf_ram.memory[135][0] ),
    .A2(_03425_),
    .ZN(_03426_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07483_ (.A1(_03306_),
    .A2(_03425_),
    .B(_03426_),
    .ZN(_00637_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07484_ (.A1(\u_cpu.rf_ram.memory[135][1] ),
    .A2(_03425_),
    .ZN(_03427_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07485_ (.A1(_03310_),
    .A2(_03425_),
    .B(_03427_),
    .ZN(_00638_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07486_ (.A1(\u_cpu.rf_ram.memory[135][2] ),
    .A2(_03425_),
    .ZN(_03428_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07487_ (.A1(_03312_),
    .A2(_03425_),
    .B(_03428_),
    .ZN(_00639_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07488_ (.A1(\u_cpu.rf_ram.memory[135][3] ),
    .A2(_03425_),
    .ZN(_03429_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07489_ (.A1(_03314_),
    .A2(_03425_),
    .B(_03429_),
    .ZN(_00640_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07490_ (.A1(\u_cpu.rf_ram.memory[135][4] ),
    .A2(_03425_),
    .ZN(_03430_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07491_ (.A1(_03316_),
    .A2(_03425_),
    .B(_03430_),
    .ZN(_00641_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07492_ (.A1(\u_cpu.rf_ram.memory[135][5] ),
    .A2(_03425_),
    .ZN(_03431_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07493_ (.A1(_03318_),
    .A2(_03425_),
    .B(_03431_),
    .ZN(_00642_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07494_ (.A1(\u_cpu.rf_ram.memory[135][6] ),
    .A2(_03425_),
    .ZN(_03432_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07495_ (.A1(_03320_),
    .A2(_03425_),
    .B(_03432_),
    .ZN(_00643_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07496_ (.A1(\u_cpu.rf_ram.memory[135][7] ),
    .A2(_03425_),
    .ZN(_03433_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07497_ (.A1(_03322_),
    .A2(_03425_),
    .B(_03433_),
    .ZN(_00644_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07498_ (.A1(_02976_),
    .A2(_03037_),
    .ZN(_03434_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07499_ (.I(_03434_),
    .Z(_03435_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07500_ (.A1(\u_cpu.rf_ram.memory[134][0] ),
    .A2(_03435_),
    .ZN(_03436_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07501_ (.A1(_03306_),
    .A2(_03435_),
    .B(_03436_),
    .ZN(_00645_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07502_ (.A1(\u_cpu.rf_ram.memory[134][1] ),
    .A2(_03435_),
    .ZN(_03437_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07503_ (.A1(_03310_),
    .A2(_03435_),
    .B(_03437_),
    .ZN(_00646_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07504_ (.A1(\u_cpu.rf_ram.memory[134][2] ),
    .A2(_03435_),
    .ZN(_03438_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07505_ (.A1(_03312_),
    .A2(_03435_),
    .B(_03438_),
    .ZN(_00647_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07506_ (.A1(\u_cpu.rf_ram.memory[134][3] ),
    .A2(_03435_),
    .ZN(_03439_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07507_ (.A1(_03314_),
    .A2(_03435_),
    .B(_03439_),
    .ZN(_00648_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07508_ (.A1(\u_cpu.rf_ram.memory[134][4] ),
    .A2(_03435_),
    .ZN(_03440_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07509_ (.A1(_03316_),
    .A2(_03435_),
    .B(_03440_),
    .ZN(_00649_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07510_ (.A1(\u_cpu.rf_ram.memory[134][5] ),
    .A2(_03435_),
    .ZN(_03441_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07511_ (.A1(_03318_),
    .A2(_03435_),
    .B(_03441_),
    .ZN(_00650_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07512_ (.A1(\u_cpu.rf_ram.memory[134][6] ),
    .A2(_03435_),
    .ZN(_03442_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07513_ (.A1(_03320_),
    .A2(_03435_),
    .B(_03442_),
    .ZN(_00651_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07514_ (.A1(\u_cpu.rf_ram.memory[134][7] ),
    .A2(_03435_),
    .ZN(_03443_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07515_ (.A1(_03322_),
    .A2(_03435_),
    .B(_03443_),
    .ZN(_00652_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07516_ (.A1(_02675_),
    .A2(_02976_),
    .ZN(_03444_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07517_ (.I(_03444_),
    .Z(_03445_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07518_ (.A1(\u_cpu.rf_ram.memory[133][0] ),
    .A2(_03445_),
    .ZN(_03446_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07519_ (.A1(_03306_),
    .A2(_03445_),
    .B(_03446_),
    .ZN(_00653_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07520_ (.A1(\u_cpu.rf_ram.memory[133][1] ),
    .A2(_03445_),
    .ZN(_03447_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07521_ (.A1(_03310_),
    .A2(_03445_),
    .B(_03447_),
    .ZN(_00654_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07522_ (.A1(\u_cpu.rf_ram.memory[133][2] ),
    .A2(_03445_),
    .ZN(_03448_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07523_ (.A1(_03312_),
    .A2(_03445_),
    .B(_03448_),
    .ZN(_00655_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07524_ (.A1(\u_cpu.rf_ram.memory[133][3] ),
    .A2(_03445_),
    .ZN(_03449_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07525_ (.A1(_03314_),
    .A2(_03445_),
    .B(_03449_),
    .ZN(_00656_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07526_ (.A1(\u_cpu.rf_ram.memory[133][4] ),
    .A2(_03445_),
    .ZN(_03450_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07527_ (.A1(_03316_),
    .A2(_03445_),
    .B(_03450_),
    .ZN(_00657_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07528_ (.A1(\u_cpu.rf_ram.memory[133][5] ),
    .A2(_03445_),
    .ZN(_03451_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07529_ (.A1(_03318_),
    .A2(_03445_),
    .B(_03451_),
    .ZN(_00658_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07530_ (.A1(\u_cpu.rf_ram.memory[133][6] ),
    .A2(_03445_),
    .ZN(_03452_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07531_ (.A1(_03320_),
    .A2(_03445_),
    .B(_03452_),
    .ZN(_00659_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07532_ (.A1(\u_cpu.rf_ram.memory[133][7] ),
    .A2(_03445_),
    .ZN(_03453_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07533_ (.A1(_03322_),
    .A2(_03445_),
    .B(_03453_),
    .ZN(_00660_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07534_ (.A1(_02717_),
    .A2(_02976_),
    .ZN(_03454_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07535_ (.I(_03454_),
    .Z(_03455_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07536_ (.A1(\u_cpu.rf_ram.memory[132][0] ),
    .A2(_03455_),
    .ZN(_03456_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07537_ (.A1(_03306_),
    .A2(_03455_),
    .B(_03456_),
    .ZN(_00661_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07538_ (.A1(\u_cpu.rf_ram.memory[132][1] ),
    .A2(_03455_),
    .ZN(_03457_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07539_ (.A1(_03310_),
    .A2(_03455_),
    .B(_03457_),
    .ZN(_00662_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07540_ (.A1(\u_cpu.rf_ram.memory[132][2] ),
    .A2(_03455_),
    .ZN(_03458_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07541_ (.A1(_03312_),
    .A2(_03455_),
    .B(_03458_),
    .ZN(_00663_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07542_ (.A1(\u_cpu.rf_ram.memory[132][3] ),
    .A2(_03455_),
    .ZN(_03459_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07543_ (.A1(_03314_),
    .A2(_03455_),
    .B(_03459_),
    .ZN(_00664_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07544_ (.A1(\u_cpu.rf_ram.memory[132][4] ),
    .A2(_03455_),
    .ZN(_03460_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07545_ (.A1(_03316_),
    .A2(_03455_),
    .B(_03460_),
    .ZN(_00665_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07546_ (.A1(\u_cpu.rf_ram.memory[132][5] ),
    .A2(_03455_),
    .ZN(_03461_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07547_ (.A1(_03318_),
    .A2(_03455_),
    .B(_03461_),
    .ZN(_00666_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07548_ (.A1(\u_cpu.rf_ram.memory[132][6] ),
    .A2(_03455_),
    .ZN(_03462_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07549_ (.A1(_03320_),
    .A2(_03455_),
    .B(_03462_),
    .ZN(_00667_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07550_ (.A1(\u_cpu.rf_ram.memory[132][7] ),
    .A2(_03455_),
    .ZN(_03463_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07551_ (.A1(_03322_),
    .A2(_03455_),
    .B(_03463_),
    .ZN(_00668_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07552_ (.A1(_02825_),
    .A2(_02976_),
    .ZN(_03464_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07553_ (.I(_03464_),
    .Z(_03465_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07554_ (.A1(\u_cpu.rf_ram.memory[131][0] ),
    .A2(_03465_),
    .ZN(_03466_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07555_ (.A1(_03306_),
    .A2(_03465_),
    .B(_03466_),
    .ZN(_00669_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07556_ (.A1(\u_cpu.rf_ram.memory[131][1] ),
    .A2(_03465_),
    .ZN(_03467_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07557_ (.A1(_03310_),
    .A2(_03465_),
    .B(_03467_),
    .ZN(_00670_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07558_ (.A1(\u_cpu.rf_ram.memory[131][2] ),
    .A2(_03465_),
    .ZN(_03468_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07559_ (.A1(_03312_),
    .A2(_03465_),
    .B(_03468_),
    .ZN(_00671_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07560_ (.A1(\u_cpu.rf_ram.memory[131][3] ),
    .A2(_03465_),
    .ZN(_03469_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07561_ (.A1(_03314_),
    .A2(_03465_),
    .B(_03469_),
    .ZN(_00672_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07562_ (.A1(\u_cpu.rf_ram.memory[131][4] ),
    .A2(_03465_),
    .ZN(_03470_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07563_ (.A1(_03316_),
    .A2(_03465_),
    .B(_03470_),
    .ZN(_00673_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07564_ (.A1(\u_cpu.rf_ram.memory[131][5] ),
    .A2(_03465_),
    .ZN(_03471_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07565_ (.A1(_03318_),
    .A2(_03465_),
    .B(_03471_),
    .ZN(_00674_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07566_ (.A1(\u_cpu.rf_ram.memory[131][6] ),
    .A2(_03465_),
    .ZN(_03472_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07567_ (.A1(_03320_),
    .A2(_03465_),
    .B(_03472_),
    .ZN(_00675_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07568_ (.A1(\u_cpu.rf_ram.memory[131][7] ),
    .A2(_03465_),
    .ZN(_03473_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07569_ (.A1(_03322_),
    .A2(_03465_),
    .B(_03473_),
    .ZN(_00676_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07570_ (.A1(_02619_),
    .A2(_02976_),
    .ZN(_03474_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07571_ (.I(_03474_),
    .Z(_03475_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07572_ (.A1(\u_cpu.rf_ram.memory[130][0] ),
    .A2(_03475_),
    .ZN(_03476_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07573_ (.A1(_03306_),
    .A2(_03475_),
    .B(_03476_),
    .ZN(_00677_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07574_ (.A1(\u_cpu.rf_ram.memory[130][1] ),
    .A2(_03475_),
    .ZN(_03477_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07575_ (.A1(_03310_),
    .A2(_03475_),
    .B(_03477_),
    .ZN(_00678_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07576_ (.A1(\u_cpu.rf_ram.memory[130][2] ),
    .A2(_03475_),
    .ZN(_03478_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07577_ (.A1(_03312_),
    .A2(_03475_),
    .B(_03478_),
    .ZN(_00679_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07578_ (.A1(\u_cpu.rf_ram.memory[130][3] ),
    .A2(_03475_),
    .ZN(_03479_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07579_ (.A1(_03314_),
    .A2(_03475_),
    .B(_03479_),
    .ZN(_00680_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07580_ (.A1(\u_cpu.rf_ram.memory[130][4] ),
    .A2(_03475_),
    .ZN(_03480_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07581_ (.A1(_03316_),
    .A2(_03475_),
    .B(_03480_),
    .ZN(_00681_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07582_ (.A1(\u_cpu.rf_ram.memory[130][5] ),
    .A2(_03475_),
    .ZN(_03481_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07583_ (.A1(_03318_),
    .A2(_03475_),
    .B(_03481_),
    .ZN(_00682_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07584_ (.A1(\u_cpu.rf_ram.memory[130][6] ),
    .A2(_03475_),
    .ZN(_03482_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07585_ (.A1(_03320_),
    .A2(_03475_),
    .B(_03482_),
    .ZN(_00683_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07586_ (.A1(\u_cpu.rf_ram.memory[130][7] ),
    .A2(_03475_),
    .ZN(_03483_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07587_ (.A1(_03322_),
    .A2(_03475_),
    .B(_03483_),
    .ZN(_00684_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07588_ (.A1(_02731_),
    .A2(_02814_),
    .ZN(_03484_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07589_ (.I(_03484_),
    .ZN(_03485_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07590_ (.A1(\u_cpu.rf_ram.memory[12][0] ),
    .A2(_03485_),
    .ZN(_03486_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07591_ (.A1(_02632_),
    .A2(_03485_),
    .B(_03486_),
    .ZN(_00685_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07592_ (.A1(\u_cpu.rf_ram.memory[12][1] ),
    .A2(_03485_),
    .ZN(_03487_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07593_ (.A1(_02637_),
    .A2(_03485_),
    .B(_03487_),
    .ZN(_00686_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07594_ (.A1(\u_cpu.rf_ram.memory[12][2] ),
    .A2(_03485_),
    .ZN(_03488_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07595_ (.A1(_02642_),
    .A2(_03485_),
    .B(_03488_),
    .ZN(_00687_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07596_ (.A1(\u_cpu.rf_ram.memory[12][3] ),
    .A2(_03485_),
    .ZN(_03489_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07597_ (.A1(_02647_),
    .A2(_03485_),
    .B(_03489_),
    .ZN(_00688_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07598_ (.A1(\u_cpu.rf_ram.memory[12][4] ),
    .A2(_03485_),
    .ZN(_03490_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07599_ (.A1(_02652_),
    .A2(_03485_),
    .B(_03490_),
    .ZN(_00689_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07600_ (.A1(\u_cpu.rf_ram.memory[12][5] ),
    .A2(_03485_),
    .ZN(_03491_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07601_ (.A1(_02657_),
    .A2(_03485_),
    .B(_03491_),
    .ZN(_00690_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07602_ (.A1(\u_cpu.rf_ram.memory[12][6] ),
    .A2(_03485_),
    .ZN(_03492_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07603_ (.A1(_02662_),
    .A2(_03485_),
    .B(_03492_),
    .ZN(_00691_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07604_ (.A1(\u_cpu.rf_ram.memory[12][7] ),
    .A2(_03485_),
    .ZN(_03493_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07605_ (.A1(_02667_),
    .A2(_03485_),
    .B(_03493_),
    .ZN(_00692_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07606_ (.I(_02631_),
    .Z(_03494_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07607_ (.A1(_02677_),
    .A2(_03037_),
    .ZN(_03495_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07608_ (.I(_03495_),
    .Z(_03496_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07609_ (.A1(\u_cpu.rf_ram.memory[22][0] ),
    .A2(_03496_),
    .ZN(_03497_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07610_ (.A1(_03494_),
    .A2(_03496_),
    .B(_03497_),
    .ZN(_00693_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07611_ (.I(_02636_),
    .Z(_03498_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07612_ (.A1(\u_cpu.rf_ram.memory[22][1] ),
    .A2(_03496_),
    .ZN(_03499_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07613_ (.A1(_03498_),
    .A2(_03496_),
    .B(_03499_),
    .ZN(_00694_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07614_ (.I(_02641_),
    .Z(_03500_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07615_ (.A1(\u_cpu.rf_ram.memory[22][2] ),
    .A2(_03496_),
    .ZN(_03501_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07616_ (.A1(_03500_),
    .A2(_03496_),
    .B(_03501_),
    .ZN(_00695_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07617_ (.I(_02646_),
    .Z(_03502_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07618_ (.A1(\u_cpu.rf_ram.memory[22][3] ),
    .A2(_03496_),
    .ZN(_03503_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07619_ (.A1(_03502_),
    .A2(_03496_),
    .B(_03503_),
    .ZN(_00696_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07620_ (.I(_02651_),
    .Z(_03504_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07621_ (.A1(\u_cpu.rf_ram.memory[22][4] ),
    .A2(_03496_),
    .ZN(_03505_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07622_ (.A1(_03504_),
    .A2(_03496_),
    .B(_03505_),
    .ZN(_00697_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07623_ (.I(_02656_),
    .Z(_03506_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07624_ (.A1(\u_cpu.rf_ram.memory[22][5] ),
    .A2(_03496_),
    .ZN(_03507_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07625_ (.A1(_03506_),
    .A2(_03496_),
    .B(_03507_),
    .ZN(_00698_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07626_ (.I(_02661_),
    .Z(_03508_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07627_ (.A1(\u_cpu.rf_ram.memory[22][6] ),
    .A2(_03496_),
    .ZN(_03509_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07628_ (.A1(_03508_),
    .A2(_03496_),
    .B(_03509_),
    .ZN(_00699_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07629_ (.I(_02666_),
    .Z(_03510_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07630_ (.A1(\u_cpu.rf_ram.memory[22][7] ),
    .A2(_03496_),
    .ZN(_03511_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07631_ (.A1(_03510_),
    .A2(_03496_),
    .B(_03511_),
    .ZN(_00700_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07632_ (.A1(_02754_),
    .A2(_02976_),
    .ZN(_03512_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07633_ (.I(_03512_),
    .Z(_03513_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07634_ (.A1(\u_cpu.rf_ram.memory[128][0] ),
    .A2(_03513_),
    .ZN(_03514_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07635_ (.A1(_03494_),
    .A2(_03513_),
    .B(_03514_),
    .ZN(_00701_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07636_ (.A1(\u_cpu.rf_ram.memory[128][1] ),
    .A2(_03513_),
    .ZN(_03515_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07637_ (.A1(_03498_),
    .A2(_03513_),
    .B(_03515_),
    .ZN(_00702_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07638_ (.A1(\u_cpu.rf_ram.memory[128][2] ),
    .A2(_03513_),
    .ZN(_03516_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07639_ (.A1(_03500_),
    .A2(_03513_),
    .B(_03516_),
    .ZN(_00703_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07640_ (.A1(\u_cpu.rf_ram.memory[128][3] ),
    .A2(_03513_),
    .ZN(_03517_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07641_ (.A1(_03502_),
    .A2(_03513_),
    .B(_03517_),
    .ZN(_00704_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07642_ (.A1(\u_cpu.rf_ram.memory[128][4] ),
    .A2(_03513_),
    .ZN(_03518_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07643_ (.A1(_03504_),
    .A2(_03513_),
    .B(_03518_),
    .ZN(_00705_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07644_ (.A1(\u_cpu.rf_ram.memory[128][5] ),
    .A2(_03513_),
    .ZN(_03519_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07645_ (.A1(_03506_),
    .A2(_03513_),
    .B(_03519_),
    .ZN(_00706_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07646_ (.A1(\u_cpu.rf_ram.memory[128][6] ),
    .A2(_03513_),
    .ZN(_03520_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07647_ (.A1(_03508_),
    .A2(_03513_),
    .B(_03520_),
    .ZN(_00707_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07648_ (.A1(\u_cpu.rf_ram.memory[128][7] ),
    .A2(_03513_),
    .ZN(_03521_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07649_ (.A1(_03510_),
    .A2(_03513_),
    .B(_03521_),
    .ZN(_00708_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07650_ (.A1(_02870_),
    .A2(_02965_),
    .ZN(_03522_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07651_ (.I(_03522_),
    .Z(_03523_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07652_ (.A1(\u_cpu.rf_ram.memory[127][0] ),
    .A2(_03523_),
    .ZN(_03524_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07653_ (.A1(_03494_),
    .A2(_03523_),
    .B(_03524_),
    .ZN(_00709_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07654_ (.A1(\u_cpu.rf_ram.memory[127][1] ),
    .A2(_03523_),
    .ZN(_03525_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07655_ (.A1(_03498_),
    .A2(_03523_),
    .B(_03525_),
    .ZN(_00710_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07656_ (.A1(\u_cpu.rf_ram.memory[127][2] ),
    .A2(_03523_),
    .ZN(_03526_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07657_ (.A1(_03500_),
    .A2(_03523_),
    .B(_03526_),
    .ZN(_00711_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07658_ (.A1(\u_cpu.rf_ram.memory[127][3] ),
    .A2(_03523_),
    .ZN(_03527_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07659_ (.A1(_03502_),
    .A2(_03523_),
    .B(_03527_),
    .ZN(_00712_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07660_ (.A1(\u_cpu.rf_ram.memory[127][4] ),
    .A2(_03523_),
    .ZN(_03528_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07661_ (.A1(_03504_),
    .A2(_03523_),
    .B(_03528_),
    .ZN(_00713_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07662_ (.A1(\u_cpu.rf_ram.memory[127][5] ),
    .A2(_03523_),
    .ZN(_03529_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07663_ (.A1(_03506_),
    .A2(_03523_),
    .B(_03529_),
    .ZN(_00714_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07664_ (.A1(\u_cpu.rf_ram.memory[127][6] ),
    .A2(_03523_),
    .ZN(_03530_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07665_ (.A1(_03508_),
    .A2(_03523_),
    .B(_03530_),
    .ZN(_00715_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07666_ (.A1(\u_cpu.rf_ram.memory[127][7] ),
    .A2(_03523_),
    .ZN(_03531_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07667_ (.A1(_03510_),
    .A2(_03523_),
    .B(_03531_),
    .ZN(_00716_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07668_ (.A1(_02766_),
    .A2(_02965_),
    .ZN(_03532_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07669_ (.I(_03532_),
    .Z(_03533_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07670_ (.A1(\u_cpu.rf_ram.memory[126][0] ),
    .A2(_03533_),
    .ZN(_03534_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07671_ (.A1(_03494_),
    .A2(_03533_),
    .B(_03534_),
    .ZN(_00717_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07672_ (.A1(\u_cpu.rf_ram.memory[126][1] ),
    .A2(_03533_),
    .ZN(_03535_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07673_ (.A1(_03498_),
    .A2(_03533_),
    .B(_03535_),
    .ZN(_00718_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07674_ (.A1(\u_cpu.rf_ram.memory[126][2] ),
    .A2(_03533_),
    .ZN(_03536_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07675_ (.A1(_03500_),
    .A2(_03533_),
    .B(_03536_),
    .ZN(_00719_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07676_ (.A1(\u_cpu.rf_ram.memory[126][3] ),
    .A2(_03533_),
    .ZN(_03537_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07677_ (.A1(_03502_),
    .A2(_03533_),
    .B(_03537_),
    .ZN(_00720_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07678_ (.A1(\u_cpu.rf_ram.memory[126][4] ),
    .A2(_03533_),
    .ZN(_03538_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07679_ (.A1(_03504_),
    .A2(_03533_),
    .B(_03538_),
    .ZN(_00721_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07680_ (.A1(\u_cpu.rf_ram.memory[126][5] ),
    .A2(_03533_),
    .ZN(_03539_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07681_ (.A1(_03506_),
    .A2(_03533_),
    .B(_03539_),
    .ZN(_00722_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07682_ (.A1(\u_cpu.rf_ram.memory[126][6] ),
    .A2(_03533_),
    .ZN(_03540_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07683_ (.A1(_03508_),
    .A2(_03533_),
    .B(_03540_),
    .ZN(_00723_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07684_ (.A1(\u_cpu.rf_ram.memory[126][7] ),
    .A2(_03533_),
    .ZN(_03541_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07685_ (.A1(_03510_),
    .A2(_03533_),
    .B(_03541_),
    .ZN(_00724_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07686_ (.A1(_02803_),
    .A2(_02965_),
    .ZN(_03542_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07687_ (.I(_03542_),
    .Z(_03543_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07688_ (.A1(\u_cpu.rf_ram.memory[125][0] ),
    .A2(_03543_),
    .ZN(_03544_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07689_ (.A1(_03494_),
    .A2(_03543_),
    .B(_03544_),
    .ZN(_00725_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07690_ (.A1(\u_cpu.rf_ram.memory[125][1] ),
    .A2(_03543_),
    .ZN(_03545_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07691_ (.A1(_03498_),
    .A2(_03543_),
    .B(_03545_),
    .ZN(_00726_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07692_ (.A1(\u_cpu.rf_ram.memory[125][2] ),
    .A2(_03543_),
    .ZN(_03546_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07693_ (.A1(_03500_),
    .A2(_03543_),
    .B(_03546_),
    .ZN(_00727_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07694_ (.A1(\u_cpu.rf_ram.memory[125][3] ),
    .A2(_03543_),
    .ZN(_03547_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07695_ (.A1(_03502_),
    .A2(_03543_),
    .B(_03547_),
    .ZN(_00728_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07696_ (.A1(\u_cpu.rf_ram.memory[125][4] ),
    .A2(_03543_),
    .ZN(_03548_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07697_ (.A1(_03504_),
    .A2(_03543_),
    .B(_03548_),
    .ZN(_00729_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07698_ (.A1(\u_cpu.rf_ram.memory[125][5] ),
    .A2(_03543_),
    .ZN(_03549_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07699_ (.A1(_03506_),
    .A2(_03543_),
    .B(_03549_),
    .ZN(_00730_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07700_ (.A1(\u_cpu.rf_ram.memory[125][6] ),
    .A2(_03543_),
    .ZN(_03550_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07701_ (.A1(_03508_),
    .A2(_03543_),
    .B(_03550_),
    .ZN(_00731_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07702_ (.A1(\u_cpu.rf_ram.memory[125][7] ),
    .A2(_03543_),
    .ZN(_03551_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07703_ (.A1(_03510_),
    .A2(_03543_),
    .B(_03551_),
    .ZN(_00732_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07704_ (.A1(_02814_),
    .A2(_02965_),
    .ZN(_03552_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07705_ (.I(_03552_),
    .Z(_03553_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07706_ (.A1(\u_cpu.rf_ram.memory[124][0] ),
    .A2(_03553_),
    .ZN(_03554_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07707_ (.A1(_03494_),
    .A2(_03553_),
    .B(_03554_),
    .ZN(_00733_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07708_ (.A1(\u_cpu.rf_ram.memory[124][1] ),
    .A2(_03553_),
    .ZN(_03555_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07709_ (.A1(_03498_),
    .A2(_03553_),
    .B(_03555_),
    .ZN(_00734_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07710_ (.A1(\u_cpu.rf_ram.memory[124][2] ),
    .A2(_03553_),
    .ZN(_03556_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07711_ (.A1(_03500_),
    .A2(_03553_),
    .B(_03556_),
    .ZN(_00735_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07712_ (.A1(\u_cpu.rf_ram.memory[124][3] ),
    .A2(_03553_),
    .ZN(_03557_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07713_ (.A1(_03502_),
    .A2(_03553_),
    .B(_03557_),
    .ZN(_00736_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07714_ (.A1(\u_cpu.rf_ram.memory[124][4] ),
    .A2(_03553_),
    .ZN(_03558_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07715_ (.A1(_03504_),
    .A2(_03553_),
    .B(_03558_),
    .ZN(_00737_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07716_ (.A1(\u_cpu.rf_ram.memory[124][5] ),
    .A2(_03553_),
    .ZN(_03559_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07717_ (.A1(_03506_),
    .A2(_03553_),
    .B(_03559_),
    .ZN(_00738_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07718_ (.A1(\u_cpu.rf_ram.memory[124][6] ),
    .A2(_03553_),
    .ZN(_03560_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07719_ (.A1(_03508_),
    .A2(_03553_),
    .B(_03560_),
    .ZN(_00739_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07720_ (.A1(\u_cpu.rf_ram.memory[124][7] ),
    .A2(_03553_),
    .ZN(_03561_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07721_ (.A1(_03510_),
    .A2(_03553_),
    .B(_03561_),
    .ZN(_00740_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07722_ (.A1(_02849_),
    .A2(_02965_),
    .ZN(_03562_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07723_ (.I(_03562_),
    .Z(_03563_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07724_ (.A1(\u_cpu.rf_ram.memory[123][0] ),
    .A2(_03563_),
    .ZN(_03564_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07725_ (.A1(_03494_),
    .A2(_03563_),
    .B(_03564_),
    .ZN(_00741_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07726_ (.A1(\u_cpu.rf_ram.memory[123][1] ),
    .A2(_03563_),
    .ZN(_03565_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07727_ (.A1(_03498_),
    .A2(_03563_),
    .B(_03565_),
    .ZN(_00742_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07728_ (.A1(\u_cpu.rf_ram.memory[123][2] ),
    .A2(_03563_),
    .ZN(_03566_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07729_ (.A1(_03500_),
    .A2(_03563_),
    .B(_03566_),
    .ZN(_00743_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07730_ (.A1(\u_cpu.rf_ram.memory[123][3] ),
    .A2(_03563_),
    .ZN(_03567_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07731_ (.A1(_03502_),
    .A2(_03563_),
    .B(_03567_),
    .ZN(_00744_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07732_ (.A1(\u_cpu.rf_ram.memory[123][4] ),
    .A2(_03563_),
    .ZN(_03568_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07733_ (.A1(_03504_),
    .A2(_03563_),
    .B(_03568_),
    .ZN(_00745_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07734_ (.A1(\u_cpu.rf_ram.memory[123][5] ),
    .A2(_03563_),
    .ZN(_03569_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07735_ (.A1(_03506_),
    .A2(_03563_),
    .B(_03569_),
    .ZN(_00746_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07736_ (.A1(\u_cpu.rf_ram.memory[123][6] ),
    .A2(_03563_),
    .ZN(_03570_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07737_ (.A1(_03508_),
    .A2(_03563_),
    .B(_03570_),
    .ZN(_00747_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07738_ (.A1(\u_cpu.rf_ram.memory[123][7] ),
    .A2(_03563_),
    .ZN(_03571_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07739_ (.A1(_03510_),
    .A2(_03563_),
    .B(_03571_),
    .ZN(_00748_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07740_ (.A1(_02782_),
    .A2(_03037_),
    .ZN(_03572_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07741_ (.I(_03572_),
    .Z(_03573_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07742_ (.A1(\u_cpu.rf_ram.memory[38][0] ),
    .A2(_03573_),
    .ZN(_03574_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07743_ (.A1(_03494_),
    .A2(_03573_),
    .B(_03574_),
    .ZN(_00749_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07744_ (.A1(\u_cpu.rf_ram.memory[38][1] ),
    .A2(_03573_),
    .ZN(_03575_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07745_ (.A1(_03498_),
    .A2(_03573_),
    .B(_03575_),
    .ZN(_00750_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07746_ (.A1(\u_cpu.rf_ram.memory[38][2] ),
    .A2(_03573_),
    .ZN(_03576_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07747_ (.A1(_03500_),
    .A2(_03573_),
    .B(_03576_),
    .ZN(_00751_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07748_ (.A1(\u_cpu.rf_ram.memory[38][3] ),
    .A2(_03573_),
    .ZN(_03577_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07749_ (.A1(_03502_),
    .A2(_03573_),
    .B(_03577_),
    .ZN(_00752_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07750_ (.A1(\u_cpu.rf_ram.memory[38][4] ),
    .A2(_03573_),
    .ZN(_03578_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07751_ (.A1(_03504_),
    .A2(_03573_),
    .B(_03578_),
    .ZN(_00753_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07752_ (.A1(\u_cpu.rf_ram.memory[38][5] ),
    .A2(_03573_),
    .ZN(_03579_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07753_ (.A1(_03506_),
    .A2(_03573_),
    .B(_03579_),
    .ZN(_00754_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07754_ (.A1(\u_cpu.rf_ram.memory[38][6] ),
    .A2(_03573_),
    .ZN(_03580_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07755_ (.A1(_03508_),
    .A2(_03573_),
    .B(_03580_),
    .ZN(_00755_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07756_ (.A1(\u_cpu.rf_ram.memory[38][7] ),
    .A2(_03573_),
    .ZN(_03581_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07757_ (.A1(_03510_),
    .A2(_03573_),
    .B(_03581_),
    .ZN(_00756_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07758_ (.A1(_02675_),
    .A2(_02782_),
    .ZN(_03582_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07759_ (.I(_03582_),
    .Z(_03583_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07760_ (.A1(\u_cpu.rf_ram.memory[37][0] ),
    .A2(_03583_),
    .ZN(_03584_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07761_ (.A1(_03494_),
    .A2(_03583_),
    .B(_03584_),
    .ZN(_00757_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07762_ (.A1(\u_cpu.rf_ram.memory[37][1] ),
    .A2(_03583_),
    .ZN(_03585_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07763_ (.A1(_03498_),
    .A2(_03583_),
    .B(_03585_),
    .ZN(_00758_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07764_ (.A1(\u_cpu.rf_ram.memory[37][2] ),
    .A2(_03583_),
    .ZN(_03586_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07765_ (.A1(_03500_),
    .A2(_03583_),
    .B(_03586_),
    .ZN(_00759_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07766_ (.A1(\u_cpu.rf_ram.memory[37][3] ),
    .A2(_03583_),
    .ZN(_03587_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07767_ (.A1(_03502_),
    .A2(_03583_),
    .B(_03587_),
    .ZN(_00760_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07768_ (.A1(\u_cpu.rf_ram.memory[37][4] ),
    .A2(_03583_),
    .ZN(_03588_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07769_ (.A1(_03504_),
    .A2(_03583_),
    .B(_03588_),
    .ZN(_00761_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07770_ (.A1(\u_cpu.rf_ram.memory[37][5] ),
    .A2(_03583_),
    .ZN(_03589_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07771_ (.A1(_03506_),
    .A2(_03583_),
    .B(_03589_),
    .ZN(_00762_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07772_ (.A1(\u_cpu.rf_ram.memory[37][6] ),
    .A2(_03583_),
    .ZN(_03590_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07773_ (.A1(_03508_),
    .A2(_03583_),
    .B(_03590_),
    .ZN(_00763_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07774_ (.A1(\u_cpu.rf_ram.memory[37][7] ),
    .A2(_03583_),
    .ZN(_03591_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07775_ (.A1(_03510_),
    .A2(_03583_),
    .B(_03591_),
    .ZN(_00764_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07776_ (.A1(_02717_),
    .A2(_02782_),
    .ZN(_03592_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07777_ (.I(_03592_),
    .Z(_03593_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07778_ (.A1(\u_cpu.rf_ram.memory[36][0] ),
    .A2(_03593_),
    .ZN(_03594_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07779_ (.A1(_03494_),
    .A2(_03593_),
    .B(_03594_),
    .ZN(_00765_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07780_ (.A1(\u_cpu.rf_ram.memory[36][1] ),
    .A2(_03593_),
    .ZN(_03595_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07781_ (.A1(_03498_),
    .A2(_03593_),
    .B(_03595_),
    .ZN(_00766_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07782_ (.A1(\u_cpu.rf_ram.memory[36][2] ),
    .A2(_03593_),
    .ZN(_03596_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07783_ (.A1(_03500_),
    .A2(_03593_),
    .B(_03596_),
    .ZN(_00767_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07784_ (.A1(\u_cpu.rf_ram.memory[36][3] ),
    .A2(_03593_),
    .ZN(_03597_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07785_ (.A1(_03502_),
    .A2(_03593_),
    .B(_03597_),
    .ZN(_00768_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07786_ (.A1(\u_cpu.rf_ram.memory[36][4] ),
    .A2(_03593_),
    .ZN(_03598_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07787_ (.A1(_03504_),
    .A2(_03593_),
    .B(_03598_),
    .ZN(_00769_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07788_ (.A1(\u_cpu.rf_ram.memory[36][5] ),
    .A2(_03593_),
    .ZN(_03599_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07789_ (.A1(_03506_),
    .A2(_03593_),
    .B(_03599_),
    .ZN(_00770_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07790_ (.A1(\u_cpu.rf_ram.memory[36][6] ),
    .A2(_03593_),
    .ZN(_03600_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07791_ (.A1(_03508_),
    .A2(_03593_),
    .B(_03600_),
    .ZN(_00771_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07792_ (.A1(\u_cpu.rf_ram.memory[36][7] ),
    .A2(_03593_),
    .ZN(_03601_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07793_ (.A1(_03510_),
    .A2(_03593_),
    .B(_03601_),
    .ZN(_00772_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07794_ (.A1(_02263_),
    .A2(_02914_),
    .ZN(_03602_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07795_ (.A1(_02395_),
    .A2(_03602_),
    .ZN(_03603_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07796_ (.I(_03603_),
    .Z(_00773_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07797_ (.A1(\u_cpu.cpu.state.o_cnt_r[3] ),
    .A2(\u_cpu.cpu.state.o_cnt[2] ),
    .ZN(_03604_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _07798_ (.A1(\u_cpu.cpu.state.o_cnt_r[3] ),
    .A2(\u_cpu.cpu.state.o_cnt[2] ),
    .Z(_03605_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _07799_ (.A1(_02395_),
    .A2(_03604_),
    .A3(_03605_),
    .ZN(_00774_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07800_ (.A1(_02291_),
    .A2(_03605_),
    .B(_02396_),
    .ZN(_03606_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07801_ (.A1(_02291_),
    .A2(_03605_),
    .B(_03606_),
    .ZN(_00775_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07802_ (.A1(_02291_),
    .A2(_03605_),
    .ZN(_03607_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07803_ (.A1(\u_cpu.cpu.mem_bytecnt[1] ),
    .A2(_03607_),
    .Z(_03608_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07804_ (.A1(_02395_),
    .A2(_03608_),
    .ZN(_00776_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07805_ (.I(\u_cpu.rf_ram_if.rgnt ),
    .ZN(_03609_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _07806_ (.A1(_03609_),
    .A2(_02927_),
    .Z(_03610_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07807_ (.A1(_02395_),
    .A2(_02263_),
    .ZN(_03611_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07808_ (.A1(\u_cpu.cpu.state.o_cnt_r[3] ),
    .A2(_03611_),
    .ZN(_03612_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _07809_ (.A1(_02395_),
    .A2(_02259_),
    .A3(_03610_),
    .B(_03612_),
    .ZN(_00777_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _07810_ (.A1(_02396_),
    .A2(\u_cpu.cpu.state.o_cnt_r[0] ),
    .Z(_03613_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07811_ (.I(_03613_),
    .Z(_00778_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07812_ (.A1(_02395_),
    .A2(_02359_),
    .ZN(_00779_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _07813_ (.A1(_02396_),
    .A2(\u_cpu.cpu.state.o_cnt_r[2] ),
    .Z(_03614_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07814_ (.I(_03614_),
    .Z(_00780_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07815_ (.A1(_02626_),
    .A2(_02849_),
    .ZN(_03615_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07816_ (.I(_03615_),
    .Z(_03616_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07817_ (.A1(\u_cpu.rf_ram.memory[91][0] ),
    .A2(_03616_),
    .ZN(_03617_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07818_ (.A1(_03494_),
    .A2(_03616_),
    .B(_03617_),
    .ZN(_00781_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07819_ (.A1(\u_cpu.rf_ram.memory[91][1] ),
    .A2(_03616_),
    .ZN(_03618_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07820_ (.A1(_03498_),
    .A2(_03616_),
    .B(_03618_),
    .ZN(_00782_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07821_ (.A1(\u_cpu.rf_ram.memory[91][2] ),
    .A2(_03616_),
    .ZN(_03619_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07822_ (.A1(_03500_),
    .A2(_03616_),
    .B(_03619_),
    .ZN(_00783_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07823_ (.A1(\u_cpu.rf_ram.memory[91][3] ),
    .A2(_03616_),
    .ZN(_03620_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07824_ (.A1(_03502_),
    .A2(_03616_),
    .B(_03620_),
    .ZN(_00784_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07825_ (.A1(\u_cpu.rf_ram.memory[91][4] ),
    .A2(_03616_),
    .ZN(_03621_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07826_ (.A1(_03504_),
    .A2(_03616_),
    .B(_03621_),
    .ZN(_00785_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07827_ (.A1(\u_cpu.rf_ram.memory[91][5] ),
    .A2(_03616_),
    .ZN(_03622_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07828_ (.A1(_03506_),
    .A2(_03616_),
    .B(_03622_),
    .ZN(_00786_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07829_ (.A1(\u_cpu.rf_ram.memory[91][6] ),
    .A2(_03616_),
    .ZN(_03623_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07830_ (.A1(_03508_),
    .A2(_03616_),
    .B(_03623_),
    .ZN(_00787_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07831_ (.A1(\u_cpu.rf_ram.memory[91][7] ),
    .A2(_03616_),
    .ZN(_03624_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07832_ (.A1(_03510_),
    .A2(_03616_),
    .B(_03624_),
    .ZN(_00788_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07833_ (.A1(_02626_),
    .A2(_02780_),
    .ZN(_03625_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07834_ (.I(_03625_),
    .Z(_03626_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07835_ (.A1(\u_cpu.rf_ram.memory[90][0] ),
    .A2(_03626_),
    .ZN(_03627_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07836_ (.A1(_03494_),
    .A2(_03626_),
    .B(_03627_),
    .ZN(_00789_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07837_ (.A1(\u_cpu.rf_ram.memory[90][1] ),
    .A2(_03626_),
    .ZN(_03628_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07838_ (.A1(_03498_),
    .A2(_03626_),
    .B(_03628_),
    .ZN(_00790_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07839_ (.A1(\u_cpu.rf_ram.memory[90][2] ),
    .A2(_03626_),
    .ZN(_03629_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07840_ (.A1(_03500_),
    .A2(_03626_),
    .B(_03629_),
    .ZN(_00791_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07841_ (.A1(\u_cpu.rf_ram.memory[90][3] ),
    .A2(_03626_),
    .ZN(_03630_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07842_ (.A1(_03502_),
    .A2(_03626_),
    .B(_03630_),
    .ZN(_00792_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07843_ (.A1(\u_cpu.rf_ram.memory[90][4] ),
    .A2(_03626_),
    .ZN(_03631_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07844_ (.A1(_03504_),
    .A2(_03626_),
    .B(_03631_),
    .ZN(_00793_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07845_ (.A1(\u_cpu.rf_ram.memory[90][5] ),
    .A2(_03626_),
    .ZN(_03632_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07846_ (.A1(_03506_),
    .A2(_03626_),
    .B(_03632_),
    .ZN(_00794_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07847_ (.A1(\u_cpu.rf_ram.memory[90][6] ),
    .A2(_03626_),
    .ZN(_03633_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07848_ (.A1(_03508_),
    .A2(_03626_),
    .B(_03633_),
    .ZN(_00795_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07849_ (.A1(\u_cpu.rf_ram.memory[90][7] ),
    .A2(_03626_),
    .ZN(_03634_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07850_ (.A1(_03510_),
    .A2(_03626_),
    .B(_03634_),
    .ZN(_00796_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _07851_ (.A1(_01444_),
    .A2(_02305_),
    .A3(_02391_),
    .Z(_03635_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07852_ (.A1(\u_cpu.cpu.state.genblk1.misalign_trap_sync_r ),
    .A2(_03611_),
    .ZN(_03636_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _07853_ (.A1(_02395_),
    .A2(_03602_),
    .A3(_03635_),
    .B(_03636_),
    .ZN(_00797_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07854_ (.A1(\u_cpu.cpu.ctrl.i_jump ),
    .A2(_03611_),
    .ZN(_03637_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07855_ (.A1(\u_cpu.cpu.bne_or_bge ),
    .A2(_01442_),
    .B(_01441_),
    .ZN(_03638_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07856_ (.A1(\u_cpu.cpu.alu.i_rs1 ),
    .A2(_03638_),
    .ZN(_03639_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07857_ (.A1(_02277_),
    .A2(_03638_),
    .ZN(_03640_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _07858_ (.A1(_02280_),
    .A2(_03640_),
    .ZN(_03641_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _07859_ (.A1(_03639_),
    .A2(_03641_),
    .Z(_03642_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07860_ (.A1(_02285_),
    .A2(_02309_),
    .B1(_03639_),
    .B2(_03641_),
    .ZN(_03643_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07861_ (.I(\u_cpu.cpu.alu.cmp_r ),
    .ZN(_03644_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _07862_ (.A1(_03644_),
    .A2(_02334_),
    .B(_01441_),
    .C(_01442_),
    .ZN(_03645_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07863_ (.A1(_03642_),
    .A2(_03643_),
    .B1(_03645_),
    .B2(_02348_),
    .ZN(_03646_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07864_ (.A1(_02286_),
    .A2(_03646_),
    .Z(_03647_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07865_ (.A1(_02265_),
    .A2(_03647_),
    .B(_00773_),
    .C(_02305_),
    .ZN(_03648_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07866_ (.A1(_03637_),
    .A2(_03648_),
    .ZN(_00799_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _07867_ (.A1(\u_cpu.cpu.mem_bytecnt[1] ),
    .A2(\u_cpu.cpu.state.o_cnt[2] ),
    .A3(_02291_),
    .A4(_00780_),
    .Z(_03649_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07868_ (.I(_03649_),
    .Z(_00800_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07869_ (.A1(\u_cpu.cpu.state.init_done ),
    .A2(_03611_),
    .ZN(_03650_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07870_ (.A1(_02395_),
    .A2(_03602_),
    .B(_03650_),
    .ZN(_00801_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07871_ (.A1(_02626_),
    .A2(_02814_),
    .ZN(_03651_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07872_ (.I(_03651_),
    .Z(_03652_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07873_ (.A1(\u_cpu.rf_ram.memory[92][0] ),
    .A2(_03652_),
    .ZN(_03653_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07874_ (.A1(_03494_),
    .A2(_03652_),
    .B(_03653_),
    .ZN(_00802_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07875_ (.A1(\u_cpu.rf_ram.memory[92][1] ),
    .A2(_03652_),
    .ZN(_03654_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07876_ (.A1(_03498_),
    .A2(_03652_),
    .B(_03654_),
    .ZN(_00803_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07877_ (.A1(\u_cpu.rf_ram.memory[92][2] ),
    .A2(_03652_),
    .ZN(_03655_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07878_ (.A1(_03500_),
    .A2(_03652_),
    .B(_03655_),
    .ZN(_00804_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07879_ (.A1(\u_cpu.rf_ram.memory[92][3] ),
    .A2(_03652_),
    .ZN(_03656_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07880_ (.A1(_03502_),
    .A2(_03652_),
    .B(_03656_),
    .ZN(_00805_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07881_ (.A1(\u_cpu.rf_ram.memory[92][4] ),
    .A2(_03652_),
    .ZN(_03657_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07882_ (.A1(_03504_),
    .A2(_03652_),
    .B(_03657_),
    .ZN(_00806_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07883_ (.A1(\u_cpu.rf_ram.memory[92][5] ),
    .A2(_03652_),
    .ZN(_03658_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07884_ (.A1(_03506_),
    .A2(_03652_),
    .B(_03658_),
    .ZN(_00807_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07885_ (.A1(\u_cpu.rf_ram.memory[92][6] ),
    .A2(_03652_),
    .ZN(_03659_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07886_ (.A1(_03508_),
    .A2(_03652_),
    .B(_03659_),
    .ZN(_00808_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07887_ (.A1(\u_cpu.rf_ram.memory[92][7] ),
    .A2(_03652_),
    .ZN(_03660_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07888_ (.A1(_03510_),
    .A2(_03652_),
    .B(_03660_),
    .ZN(_00809_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07889_ (.A1(_02782_),
    .A2(_02825_),
    .ZN(_03661_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07890_ (.I(_03661_),
    .Z(_03662_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07891_ (.A1(\u_cpu.rf_ram.memory[35][0] ),
    .A2(_03662_),
    .ZN(_03663_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07892_ (.A1(_03494_),
    .A2(_03662_),
    .B(_03663_),
    .ZN(_00810_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07893_ (.A1(\u_cpu.rf_ram.memory[35][1] ),
    .A2(_03662_),
    .ZN(_03664_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07894_ (.A1(_03498_),
    .A2(_03662_),
    .B(_03664_),
    .ZN(_00811_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07895_ (.A1(\u_cpu.rf_ram.memory[35][2] ),
    .A2(_03662_),
    .ZN(_03665_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07896_ (.A1(_03500_),
    .A2(_03662_),
    .B(_03665_),
    .ZN(_00812_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07897_ (.A1(\u_cpu.rf_ram.memory[35][3] ),
    .A2(_03662_),
    .ZN(_03666_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07898_ (.A1(_03502_),
    .A2(_03662_),
    .B(_03666_),
    .ZN(_00813_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07899_ (.A1(\u_cpu.rf_ram.memory[35][4] ),
    .A2(_03662_),
    .ZN(_03667_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07900_ (.A1(_03504_),
    .A2(_03662_),
    .B(_03667_),
    .ZN(_00814_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07901_ (.A1(\u_cpu.rf_ram.memory[35][5] ),
    .A2(_03662_),
    .ZN(_03668_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07902_ (.A1(_03506_),
    .A2(_03662_),
    .B(_03668_),
    .ZN(_00815_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07903_ (.A1(\u_cpu.rf_ram.memory[35][6] ),
    .A2(_03662_),
    .ZN(_03669_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07904_ (.A1(_03508_),
    .A2(_03662_),
    .B(_03669_),
    .ZN(_00816_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07905_ (.A1(\u_cpu.rf_ram.memory[35][7] ),
    .A2(_03662_),
    .ZN(_03670_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07906_ (.A1(_03510_),
    .A2(_03662_),
    .B(_03670_),
    .ZN(_00817_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07907_ (.A1(_02619_),
    .A2(_02782_),
    .ZN(_03671_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07908_ (.I(_03671_),
    .Z(_03672_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07909_ (.A1(\u_cpu.rf_ram.memory[34][0] ),
    .A2(_03672_),
    .ZN(_03673_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07910_ (.A1(_03494_),
    .A2(_03672_),
    .B(_03673_),
    .ZN(_00818_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07911_ (.A1(\u_cpu.rf_ram.memory[34][1] ),
    .A2(_03672_),
    .ZN(_03674_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07912_ (.A1(_03498_),
    .A2(_03672_),
    .B(_03674_),
    .ZN(_00819_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07913_ (.A1(\u_cpu.rf_ram.memory[34][2] ),
    .A2(_03672_),
    .ZN(_03675_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07914_ (.A1(_03500_),
    .A2(_03672_),
    .B(_03675_),
    .ZN(_00820_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07915_ (.A1(\u_cpu.rf_ram.memory[34][3] ),
    .A2(_03672_),
    .ZN(_03676_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07916_ (.A1(_03502_),
    .A2(_03672_),
    .B(_03676_),
    .ZN(_00821_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07917_ (.A1(\u_cpu.rf_ram.memory[34][4] ),
    .A2(_03672_),
    .ZN(_03677_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07918_ (.A1(_03504_),
    .A2(_03672_),
    .B(_03677_),
    .ZN(_00822_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07919_ (.A1(\u_cpu.rf_ram.memory[34][5] ),
    .A2(_03672_),
    .ZN(_03678_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07920_ (.A1(_03506_),
    .A2(_03672_),
    .B(_03678_),
    .ZN(_00823_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07921_ (.A1(\u_cpu.rf_ram.memory[34][6] ),
    .A2(_03672_),
    .ZN(_03679_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07922_ (.A1(_03508_),
    .A2(_03672_),
    .B(_03679_),
    .ZN(_00824_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07923_ (.A1(\u_cpu.rf_ram.memory[34][7] ),
    .A2(_03672_),
    .ZN(_03680_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07924_ (.A1(_03510_),
    .A2(_03672_),
    .B(_03680_),
    .ZN(_00825_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07925_ (.A1(_02675_),
    .A2(_02965_),
    .ZN(_03681_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07926_ (.I(_03681_),
    .Z(_03682_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07927_ (.A1(\u_cpu.rf_ram.memory[117][0] ),
    .A2(_03682_),
    .ZN(_03683_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07928_ (.A1(_03494_),
    .A2(_03682_),
    .B(_03683_),
    .ZN(_00826_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07929_ (.A1(\u_cpu.rf_ram.memory[117][1] ),
    .A2(_03682_),
    .ZN(_03684_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07930_ (.A1(_03498_),
    .A2(_03682_),
    .B(_03684_),
    .ZN(_00827_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07931_ (.A1(\u_cpu.rf_ram.memory[117][2] ),
    .A2(_03682_),
    .ZN(_03685_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07932_ (.A1(_03500_),
    .A2(_03682_),
    .B(_03685_),
    .ZN(_00828_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07933_ (.A1(\u_cpu.rf_ram.memory[117][3] ),
    .A2(_03682_),
    .ZN(_03686_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07934_ (.A1(_03502_),
    .A2(_03682_),
    .B(_03686_),
    .ZN(_00829_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07935_ (.A1(\u_cpu.rf_ram.memory[117][4] ),
    .A2(_03682_),
    .ZN(_03687_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07936_ (.A1(_03504_),
    .A2(_03682_),
    .B(_03687_),
    .ZN(_00830_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07937_ (.A1(\u_cpu.rf_ram.memory[117][5] ),
    .A2(_03682_),
    .ZN(_03688_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07938_ (.A1(_03506_),
    .A2(_03682_),
    .B(_03688_),
    .ZN(_00831_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07939_ (.A1(\u_cpu.rf_ram.memory[117][6] ),
    .A2(_03682_),
    .ZN(_03689_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07940_ (.A1(_03508_),
    .A2(_03682_),
    .B(_03689_),
    .ZN(_00832_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07941_ (.A1(\u_cpu.rf_ram.memory[117][7] ),
    .A2(_03682_),
    .ZN(_03690_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07942_ (.A1(_03510_),
    .A2(_03682_),
    .B(_03690_),
    .ZN(_00833_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07943_ (.I(_02631_),
    .Z(_03691_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07944_ (.A1(_02954_),
    .A2(_02965_),
    .ZN(_03692_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07945_ (.I(_03692_),
    .Z(_03693_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07946_ (.A1(\u_cpu.rf_ram.memory[120][0] ),
    .A2(_03693_),
    .ZN(_03694_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07947_ (.A1(_03691_),
    .A2(_03693_),
    .B(_03694_),
    .ZN(_00834_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07948_ (.I(_02636_),
    .Z(_03695_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07949_ (.A1(\u_cpu.rf_ram.memory[120][1] ),
    .A2(_03693_),
    .ZN(_03696_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07950_ (.A1(_03695_),
    .A2(_03693_),
    .B(_03696_),
    .ZN(_00835_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07951_ (.I(_02641_),
    .Z(_03697_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07952_ (.A1(\u_cpu.rf_ram.memory[120][2] ),
    .A2(_03693_),
    .ZN(_03698_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07953_ (.A1(_03697_),
    .A2(_03693_),
    .B(_03698_),
    .ZN(_00836_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07954_ (.I(_02646_),
    .Z(_03699_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07955_ (.A1(\u_cpu.rf_ram.memory[120][3] ),
    .A2(_03693_),
    .ZN(_03700_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07956_ (.A1(_03699_),
    .A2(_03693_),
    .B(_03700_),
    .ZN(_00837_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07957_ (.I(_02651_),
    .Z(_03701_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07958_ (.A1(\u_cpu.rf_ram.memory[120][4] ),
    .A2(_03693_),
    .ZN(_03702_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07959_ (.A1(_03701_),
    .A2(_03693_),
    .B(_03702_),
    .ZN(_00838_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07960_ (.I(_02656_),
    .Z(_03703_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07961_ (.A1(\u_cpu.rf_ram.memory[120][5] ),
    .A2(_03693_),
    .ZN(_03704_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07962_ (.A1(_03703_),
    .A2(_03693_),
    .B(_03704_),
    .ZN(_00839_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07963_ (.I(_02661_),
    .Z(_03705_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07964_ (.A1(\u_cpu.rf_ram.memory[120][6] ),
    .A2(_03693_),
    .ZN(_03706_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07965_ (.A1(_03705_),
    .A2(_03693_),
    .B(_03706_),
    .ZN(_00840_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07966_ (.I(_02666_),
    .Z(_03707_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07967_ (.A1(\u_cpu.rf_ram.memory[120][7] ),
    .A2(_03693_),
    .ZN(_03708_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07968_ (.A1(_03707_),
    .A2(_03693_),
    .B(_03708_),
    .ZN(_00841_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07969_ (.A1(_02965_),
    .A2(_03037_),
    .ZN(_03709_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07970_ (.I(_03709_),
    .Z(_03710_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07971_ (.A1(\u_cpu.rf_ram.memory[118][0] ),
    .A2(_03710_),
    .ZN(_03711_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07972_ (.A1(_03691_),
    .A2(_03710_),
    .B(_03711_),
    .ZN(_00842_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07973_ (.A1(\u_cpu.rf_ram.memory[118][1] ),
    .A2(_03710_),
    .ZN(_03712_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07974_ (.A1(_03695_),
    .A2(_03710_),
    .B(_03712_),
    .ZN(_00843_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07975_ (.A1(\u_cpu.rf_ram.memory[118][2] ),
    .A2(_03710_),
    .ZN(_03713_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07976_ (.A1(_03697_),
    .A2(_03710_),
    .B(_03713_),
    .ZN(_00844_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07977_ (.A1(\u_cpu.rf_ram.memory[118][3] ),
    .A2(_03710_),
    .ZN(_03714_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07978_ (.A1(_03699_),
    .A2(_03710_),
    .B(_03714_),
    .ZN(_00845_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07979_ (.A1(\u_cpu.rf_ram.memory[118][4] ),
    .A2(_03710_),
    .ZN(_03715_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07980_ (.A1(_03701_),
    .A2(_03710_),
    .B(_03715_),
    .ZN(_00846_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07981_ (.A1(\u_cpu.rf_ram.memory[118][5] ),
    .A2(_03710_),
    .ZN(_03716_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07982_ (.A1(_03703_),
    .A2(_03710_),
    .B(_03716_),
    .ZN(_00847_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07983_ (.A1(\u_cpu.rf_ram.memory[118][6] ),
    .A2(_03710_),
    .ZN(_03717_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07984_ (.A1(_03705_),
    .A2(_03710_),
    .B(_03717_),
    .ZN(_00848_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07985_ (.A1(\u_cpu.rf_ram.memory[118][7] ),
    .A2(_03710_),
    .ZN(_03718_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07986_ (.A1(_03707_),
    .A2(_03710_),
    .B(_03718_),
    .ZN(_00849_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07987_ (.A1(_02838_),
    .A2(_02965_),
    .ZN(_03719_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07988_ (.I(_03719_),
    .Z(_03720_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07989_ (.A1(\u_cpu.rf_ram.memory[121][0] ),
    .A2(_03720_),
    .ZN(_03721_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07990_ (.A1(_03691_),
    .A2(_03720_),
    .B(_03721_),
    .ZN(_00850_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07991_ (.A1(\u_cpu.rf_ram.memory[121][1] ),
    .A2(_03720_),
    .ZN(_03722_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07992_ (.A1(_03695_),
    .A2(_03720_),
    .B(_03722_),
    .ZN(_00851_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07993_ (.A1(\u_cpu.rf_ram.memory[121][2] ),
    .A2(_03720_),
    .ZN(_03723_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07994_ (.A1(_03697_),
    .A2(_03720_),
    .B(_03723_),
    .ZN(_00852_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07995_ (.A1(\u_cpu.rf_ram.memory[121][3] ),
    .A2(_03720_),
    .ZN(_03724_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07996_ (.A1(_03699_),
    .A2(_03720_),
    .B(_03724_),
    .ZN(_00853_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07997_ (.A1(\u_cpu.rf_ram.memory[121][4] ),
    .A2(_03720_),
    .ZN(_03725_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07998_ (.A1(_03701_),
    .A2(_03720_),
    .B(_03725_),
    .ZN(_00854_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07999_ (.A1(\u_cpu.rf_ram.memory[121][5] ),
    .A2(_03720_),
    .ZN(_03726_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08000_ (.A1(_03703_),
    .A2(_03720_),
    .B(_03726_),
    .ZN(_00855_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08001_ (.A1(\u_cpu.rf_ram.memory[121][6] ),
    .A2(_03720_),
    .ZN(_03727_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08002_ (.A1(_03705_),
    .A2(_03720_),
    .B(_03727_),
    .ZN(_00856_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08003_ (.A1(\u_cpu.rf_ram.memory[121][7] ),
    .A2(_03720_),
    .ZN(_03728_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08004_ (.A1(_03707_),
    .A2(_03720_),
    .B(_03728_),
    .ZN(_00857_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08005_ (.A1(_02731_),
    .A2(_02954_),
    .Z(_03729_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08006_ (.I(_03729_),
    .Z(_03730_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08007_ (.A1(\u_cpu.rf_ram.memory[8][0] ),
    .A2(_03730_),
    .ZN(_03731_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08008_ (.A1(_02632_),
    .A2(_03730_),
    .B(_03731_),
    .ZN(_00858_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08009_ (.A1(\u_cpu.rf_ram.memory[8][1] ),
    .A2(_03730_),
    .ZN(_03732_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08010_ (.A1(_02637_),
    .A2(_03730_),
    .B(_03732_),
    .ZN(_00859_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08011_ (.A1(\u_cpu.rf_ram.memory[8][2] ),
    .A2(_03730_),
    .ZN(_03733_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08012_ (.A1(_02642_),
    .A2(_03730_),
    .B(_03733_),
    .ZN(_00860_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08013_ (.A1(\u_cpu.rf_ram.memory[8][3] ),
    .A2(_03730_),
    .ZN(_03734_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08014_ (.A1(_02647_),
    .A2(_03730_),
    .B(_03734_),
    .ZN(_00861_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08015_ (.A1(\u_cpu.rf_ram.memory[8][4] ),
    .A2(_03730_),
    .ZN(_03735_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08016_ (.A1(_02652_),
    .A2(_03730_),
    .B(_03735_),
    .ZN(_00862_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08017_ (.A1(\u_cpu.rf_ram.memory[8][5] ),
    .A2(_03730_),
    .ZN(_03736_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08018_ (.A1(_02657_),
    .A2(_03730_),
    .B(_03736_),
    .ZN(_00863_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08019_ (.A1(\u_cpu.rf_ram.memory[8][6] ),
    .A2(_03730_),
    .ZN(_03737_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08020_ (.A1(_02662_),
    .A2(_03730_),
    .B(_03737_),
    .ZN(_00864_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08021_ (.A1(\u_cpu.rf_ram.memory[8][7] ),
    .A2(_03730_),
    .ZN(_03738_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08022_ (.A1(_02667_),
    .A2(_03730_),
    .B(_03738_),
    .ZN(_00865_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08023_ (.A1(_02731_),
    .A2(_02849_),
    .ZN(_03739_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08024_ (.I(_03739_),
    .ZN(_03740_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08025_ (.A1(\u_cpu.rf_ram.memory[11][0] ),
    .A2(_03740_),
    .ZN(_03741_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08026_ (.A1(_02632_),
    .A2(_03740_),
    .B(_03741_),
    .ZN(_00866_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08027_ (.A1(\u_cpu.rf_ram.memory[11][1] ),
    .A2(_03740_),
    .ZN(_03742_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08028_ (.A1(_02637_),
    .A2(_03740_),
    .B(_03742_),
    .ZN(_00867_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08029_ (.A1(\u_cpu.rf_ram.memory[11][2] ),
    .A2(_03740_),
    .ZN(_03743_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08030_ (.A1(_02642_),
    .A2(_03740_),
    .B(_03743_),
    .ZN(_00868_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08031_ (.A1(\u_cpu.rf_ram.memory[11][3] ),
    .A2(_03740_),
    .ZN(_03744_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08032_ (.A1(_02647_),
    .A2(_03740_),
    .B(_03744_),
    .ZN(_00869_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08033_ (.A1(\u_cpu.rf_ram.memory[11][4] ),
    .A2(_03740_),
    .ZN(_03745_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08034_ (.A1(_02652_),
    .A2(_03740_),
    .B(_03745_),
    .ZN(_00870_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08035_ (.A1(\u_cpu.rf_ram.memory[11][5] ),
    .A2(_03740_),
    .ZN(_03746_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08036_ (.A1(_02657_),
    .A2(_03740_),
    .B(_03746_),
    .ZN(_00871_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08037_ (.A1(\u_cpu.rf_ram.memory[11][6] ),
    .A2(_03740_),
    .ZN(_03747_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08038_ (.A1(_02662_),
    .A2(_03740_),
    .B(_03747_),
    .ZN(_00872_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08039_ (.A1(\u_cpu.rf_ram.memory[11][7] ),
    .A2(_03740_),
    .ZN(_03748_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08040_ (.A1(_02667_),
    .A2(_03740_),
    .B(_03748_),
    .ZN(_00873_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08041_ (.A1(_02754_),
    .A2(_02965_),
    .ZN(_03749_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08042_ (.I(_03749_),
    .Z(_03750_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08043_ (.A1(\u_cpu.rf_ram.memory[112][0] ),
    .A2(_03750_),
    .ZN(_03751_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08044_ (.A1(_03691_),
    .A2(_03750_),
    .B(_03751_),
    .ZN(_00874_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08045_ (.A1(\u_cpu.rf_ram.memory[112][1] ),
    .A2(_03750_),
    .ZN(_03752_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08046_ (.A1(_03695_),
    .A2(_03750_),
    .B(_03752_),
    .ZN(_00875_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08047_ (.A1(\u_cpu.rf_ram.memory[112][2] ),
    .A2(_03750_),
    .ZN(_03753_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08048_ (.A1(_03697_),
    .A2(_03750_),
    .B(_03753_),
    .ZN(_00876_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08049_ (.A1(\u_cpu.rf_ram.memory[112][3] ),
    .A2(_03750_),
    .ZN(_03754_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08050_ (.A1(_03699_),
    .A2(_03750_),
    .B(_03754_),
    .ZN(_00877_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08051_ (.A1(\u_cpu.rf_ram.memory[112][4] ),
    .A2(_03750_),
    .ZN(_03755_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08052_ (.A1(_03701_),
    .A2(_03750_),
    .B(_03755_),
    .ZN(_00878_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08053_ (.A1(\u_cpu.rf_ram.memory[112][5] ),
    .A2(_03750_),
    .ZN(_03756_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08054_ (.A1(_03703_),
    .A2(_03750_),
    .B(_03756_),
    .ZN(_00879_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08055_ (.A1(\u_cpu.rf_ram.memory[112][6] ),
    .A2(_03750_),
    .ZN(_03757_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08056_ (.A1(_03705_),
    .A2(_03750_),
    .B(_03757_),
    .ZN(_00880_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08057_ (.A1(\u_cpu.rf_ram.memory[112][7] ),
    .A2(_03750_),
    .ZN(_03758_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08058_ (.A1(_03707_),
    .A2(_03750_),
    .B(_03758_),
    .ZN(_00881_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08059_ (.A1(_02780_),
    .A2(_02965_),
    .ZN(_03759_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08060_ (.I(_03759_),
    .Z(_03760_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08061_ (.A1(\u_cpu.rf_ram.memory[122][0] ),
    .A2(_03760_),
    .ZN(_03761_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08062_ (.A1(_03691_),
    .A2(_03760_),
    .B(_03761_),
    .ZN(_00882_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08063_ (.A1(\u_cpu.rf_ram.memory[122][1] ),
    .A2(_03760_),
    .ZN(_03762_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08064_ (.A1(_03695_),
    .A2(_03760_),
    .B(_03762_),
    .ZN(_00883_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08065_ (.A1(\u_cpu.rf_ram.memory[122][2] ),
    .A2(_03760_),
    .ZN(_03763_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08066_ (.A1(_03697_),
    .A2(_03760_),
    .B(_03763_),
    .ZN(_00884_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08067_ (.A1(\u_cpu.rf_ram.memory[122][3] ),
    .A2(_03760_),
    .ZN(_03764_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08068_ (.A1(_03699_),
    .A2(_03760_),
    .B(_03764_),
    .ZN(_00885_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08069_ (.A1(\u_cpu.rf_ram.memory[122][4] ),
    .A2(_03760_),
    .ZN(_03765_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08070_ (.A1(_03701_),
    .A2(_03760_),
    .B(_03765_),
    .ZN(_00886_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08071_ (.A1(\u_cpu.rf_ram.memory[122][5] ),
    .A2(_03760_),
    .ZN(_03766_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08072_ (.A1(_03703_),
    .A2(_03760_),
    .B(_03766_),
    .ZN(_00887_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08073_ (.A1(\u_cpu.rf_ram.memory[122][6] ),
    .A2(_03760_),
    .ZN(_03767_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08074_ (.A1(_03705_),
    .A2(_03760_),
    .B(_03767_),
    .ZN(_00888_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08075_ (.A1(\u_cpu.rf_ram.memory[122][7] ),
    .A2(_03760_),
    .ZN(_03768_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08076_ (.A1(_03707_),
    .A2(_03760_),
    .B(_03768_),
    .ZN(_00889_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08077_ (.A1(_02825_),
    .A2(_02965_),
    .ZN(_03769_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08078_ (.I(_03769_),
    .Z(_03770_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08079_ (.A1(\u_cpu.rf_ram.memory[115][0] ),
    .A2(_03770_),
    .ZN(_03771_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08080_ (.A1(_03691_),
    .A2(_03770_),
    .B(_03771_),
    .ZN(_00890_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08081_ (.A1(\u_cpu.rf_ram.memory[115][1] ),
    .A2(_03770_),
    .ZN(_03772_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08082_ (.A1(_03695_),
    .A2(_03770_),
    .B(_03772_),
    .ZN(_00891_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08083_ (.A1(\u_cpu.rf_ram.memory[115][2] ),
    .A2(_03770_),
    .ZN(_03773_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08084_ (.A1(_03697_),
    .A2(_03770_),
    .B(_03773_),
    .ZN(_00892_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08085_ (.A1(\u_cpu.rf_ram.memory[115][3] ),
    .A2(_03770_),
    .ZN(_03774_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08086_ (.A1(_03699_),
    .A2(_03770_),
    .B(_03774_),
    .ZN(_00893_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08087_ (.A1(\u_cpu.rf_ram.memory[115][4] ),
    .A2(_03770_),
    .ZN(_03775_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08088_ (.A1(_03701_),
    .A2(_03770_),
    .B(_03775_),
    .ZN(_00894_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08089_ (.A1(\u_cpu.rf_ram.memory[115][5] ),
    .A2(_03770_),
    .ZN(_03776_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08090_ (.A1(_03703_),
    .A2(_03770_),
    .B(_03776_),
    .ZN(_00895_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08091_ (.A1(\u_cpu.rf_ram.memory[115][6] ),
    .A2(_03770_),
    .ZN(_03777_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08092_ (.A1(_03705_),
    .A2(_03770_),
    .B(_03777_),
    .ZN(_00896_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08093_ (.A1(\u_cpu.rf_ram.memory[115][7] ),
    .A2(_03770_),
    .ZN(_03778_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08094_ (.A1(_03707_),
    .A2(_03770_),
    .B(_03778_),
    .ZN(_00897_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08095_ (.A1(_02717_),
    .A2(_02965_),
    .ZN(_03779_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08096_ (.I(_03779_),
    .Z(_03780_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08097_ (.A1(\u_cpu.rf_ram.memory[116][0] ),
    .A2(_03780_),
    .ZN(_03781_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08098_ (.A1(_03691_),
    .A2(_03780_),
    .B(_03781_),
    .ZN(_00898_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08099_ (.A1(\u_cpu.rf_ram.memory[116][1] ),
    .A2(_03780_),
    .ZN(_03782_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08100_ (.A1(_03695_),
    .A2(_03780_),
    .B(_03782_),
    .ZN(_00899_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08101_ (.A1(\u_cpu.rf_ram.memory[116][2] ),
    .A2(_03780_),
    .ZN(_03783_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08102_ (.A1(_03697_),
    .A2(_03780_),
    .B(_03783_),
    .ZN(_00900_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08103_ (.A1(\u_cpu.rf_ram.memory[116][3] ),
    .A2(_03780_),
    .ZN(_03784_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08104_ (.A1(_03699_),
    .A2(_03780_),
    .B(_03784_),
    .ZN(_00901_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08105_ (.A1(\u_cpu.rf_ram.memory[116][4] ),
    .A2(_03780_),
    .ZN(_03785_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08106_ (.A1(_03701_),
    .A2(_03780_),
    .B(_03785_),
    .ZN(_00902_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08107_ (.A1(\u_cpu.rf_ram.memory[116][5] ),
    .A2(_03780_),
    .ZN(_03786_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08108_ (.A1(_03703_),
    .A2(_03780_),
    .B(_03786_),
    .ZN(_00903_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08109_ (.A1(\u_cpu.rf_ram.memory[116][6] ),
    .A2(_03780_),
    .ZN(_03787_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08110_ (.A1(_03705_),
    .A2(_03780_),
    .B(_03787_),
    .ZN(_00904_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08111_ (.A1(\u_cpu.rf_ram.memory[116][7] ),
    .A2(_03780_),
    .ZN(_03788_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08112_ (.A1(_03707_),
    .A2(_03780_),
    .B(_03788_),
    .ZN(_00905_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08113_ (.A1(_02695_),
    .A2(_02782_),
    .ZN(_03789_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08114_ (.I(_03789_),
    .Z(_03790_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08115_ (.A1(\u_cpu.rf_ram.memory[33][0] ),
    .A2(_03790_),
    .ZN(_03791_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08116_ (.A1(_03691_),
    .A2(_03790_),
    .B(_03791_),
    .ZN(_00906_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08117_ (.A1(\u_cpu.rf_ram.memory[33][1] ),
    .A2(_03790_),
    .ZN(_03792_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08118_ (.A1(_03695_),
    .A2(_03790_),
    .B(_03792_),
    .ZN(_00907_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08119_ (.A1(\u_cpu.rf_ram.memory[33][2] ),
    .A2(_03790_),
    .ZN(_03793_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08120_ (.A1(_03697_),
    .A2(_03790_),
    .B(_03793_),
    .ZN(_00908_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08121_ (.A1(\u_cpu.rf_ram.memory[33][3] ),
    .A2(_03790_),
    .ZN(_03794_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08122_ (.A1(_03699_),
    .A2(_03790_),
    .B(_03794_),
    .ZN(_00909_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08123_ (.A1(\u_cpu.rf_ram.memory[33][4] ),
    .A2(_03790_),
    .ZN(_03795_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08124_ (.A1(_03701_),
    .A2(_03790_),
    .B(_03795_),
    .ZN(_00910_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08125_ (.A1(\u_cpu.rf_ram.memory[33][5] ),
    .A2(_03790_),
    .ZN(_03796_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08126_ (.A1(_03703_),
    .A2(_03790_),
    .B(_03796_),
    .ZN(_00911_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08127_ (.A1(\u_cpu.rf_ram.memory[33][6] ),
    .A2(_03790_),
    .ZN(_03797_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08128_ (.A1(_03705_),
    .A2(_03790_),
    .B(_03797_),
    .ZN(_00912_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08129_ (.A1(\u_cpu.rf_ram.memory[33][7] ),
    .A2(_03790_),
    .ZN(_03798_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08130_ (.A1(_03707_),
    .A2(_03790_),
    .B(_03798_),
    .ZN(_00913_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08131_ (.A1(\u_cpu.cpu.mem_bytecnt[1] ),
    .A2(_02355_),
    .B(_02306_),
    .C(_02291_),
    .ZN(_03799_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08132_ (.A1(\u_cpu.cpu.mem_bytecnt[1] ),
    .A2(_02355_),
    .ZN(_03800_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08133_ (.A1(_02259_),
    .A2(_03799_),
    .A3(_03800_),
    .ZN(_03801_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08134_ (.A1(_02913_),
    .A2(_03801_),
    .ZN(_03802_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08135_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[0] ),
    .A2(_02915_),
    .ZN(_03803_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08136_ (.A1(_03802_),
    .A2(_03803_),
    .ZN(_03804_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08137_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[1] ),
    .A2(_02915_),
    .B(_02924_),
    .ZN(_03805_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08138_ (.A1(\u_arbiter.i_wb_cpu_ack ),
    .A2(_02397_),
    .Z(_03806_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08139_ (.I(_03806_),
    .Z(_03807_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08140_ (.A1(_03807_),
    .A2(_03802_),
    .ZN(_03808_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08141_ (.A1(\u_arbiter.i_wb_cpu_rdt[0] ),
    .A2(_03807_),
    .B1(_03808_),
    .B2(\u_arbiter.i_wb_cpu_dbus_dat[0] ),
    .ZN(_03809_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08142_ (.A1(_03804_),
    .A2(_03805_),
    .B(_03809_),
    .ZN(_00914_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08143_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[2] ),
    .A2(_02915_),
    .ZN(_03810_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08144_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[0] ),
    .A2(\u_arbiter.i_wb_cpu_dbus_dat[1] ),
    .B(_02915_),
    .ZN(_03811_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08145_ (.A1(_03802_),
    .A2(_03811_),
    .ZN(_03812_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08146_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[1] ),
    .A2(_03804_),
    .ZN(_03813_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08147_ (.A1(_03810_),
    .A2(_03812_),
    .B(_02924_),
    .C(_03813_),
    .ZN(_03814_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08148_ (.A1(\u_arbiter.i_wb_cpu_rdt[1] ),
    .A2(_02924_),
    .B(_03814_),
    .ZN(_03815_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _08149_ (.I(_03815_),
    .ZN(_00915_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08150_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[3] ),
    .A2(_02915_),
    .ZN(_03816_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _08151_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[2] ),
    .A2(\u_arbiter.i_wb_cpu_dbus_dat[0] ),
    .A3(\u_arbiter.i_wb_cpu_dbus_dat[1] ),
    .B(_02915_),
    .ZN(_03817_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08152_ (.A1(_03802_),
    .A2(_03817_),
    .ZN(_03818_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08153_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[2] ),
    .A2(_03812_),
    .ZN(_03819_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08154_ (.A1(_03816_),
    .A2(_03818_),
    .B(_02924_),
    .C(_03819_),
    .ZN(_03820_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08155_ (.A1(\u_arbiter.i_wb_cpu_rdt[2] ),
    .A2(_02924_),
    .B(_03820_),
    .ZN(_03821_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _08156_ (.I(_03821_),
    .ZN(_00916_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08157_ (.I(_03807_),
    .Z(_03822_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08158_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[4] ),
    .A2(_02915_),
    .ZN(_03823_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08159_ (.A1(_02915_),
    .A2(_02916_),
    .B(_03823_),
    .ZN(_03824_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _08160_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[3] ),
    .A2(_03818_),
    .B1(_03824_),
    .B2(_03802_),
    .C(_03807_),
    .ZN(_03825_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08161_ (.A1(_02416_),
    .A2(_03822_),
    .B(_03825_),
    .ZN(_00917_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08162_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[4] ),
    .A2(_02916_),
    .Z(_03826_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08163_ (.A1(_02915_),
    .A2(_03826_),
    .ZN(_03827_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08164_ (.A1(_02924_),
    .A2(_03802_),
    .Z(_03828_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08165_ (.I(_03828_),
    .Z(_03829_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08166_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[5] ),
    .A2(_02915_),
    .B(_03827_),
    .C(_03829_),
    .ZN(_03830_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08167_ (.A1(\u_arbiter.i_wb_cpu_rdt[4] ),
    .A2(_03822_),
    .B1(_03808_),
    .B2(\u_arbiter.i_wb_cpu_dbus_dat[4] ),
    .ZN(_03831_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08168_ (.A1(_03830_),
    .A2(_03831_),
    .ZN(_00918_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08169_ (.A1(\u_arbiter.i_wb_cpu_rdt[5] ),
    .A2(_03822_),
    .ZN(_03832_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08170_ (.I(_03829_),
    .Z(_03833_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08171_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[5] ),
    .A2(_03808_),
    .B1(_03833_),
    .B2(_02922_),
    .ZN(_03834_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08172_ (.A1(_03832_),
    .A2(_03834_),
    .ZN(_00919_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08173_ (.I(_03808_),
    .Z(_03835_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08174_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[6] ),
    .A2(_03835_),
    .ZN(_03836_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08175_ (.A1(\u_arbiter.i_wb_cpu_rdt[6] ),
    .A2(_03822_),
    .B1(_03833_),
    .B2(\u_arbiter.i_wb_cpu_dbus_dat[7] ),
    .ZN(_03837_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08176_ (.A1(_03836_),
    .A2(_03837_),
    .ZN(_00920_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08177_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[7] ),
    .A2(_03835_),
    .ZN(_03838_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08178_ (.A1(\u_arbiter.i_wb_cpu_rdt[7] ),
    .A2(_03822_),
    .B1(_03833_),
    .B2(\u_arbiter.i_wb_cpu_dbus_dat[8] ),
    .ZN(_03839_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08179_ (.A1(_03838_),
    .A2(_03839_),
    .ZN(_00921_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08180_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[8] ),
    .A2(_03835_),
    .ZN(_03840_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08181_ (.A1(\u_arbiter.i_wb_cpu_rdt[8] ),
    .A2(_03822_),
    .B1(_03833_),
    .B2(\u_arbiter.i_wb_cpu_dbus_dat[9] ),
    .ZN(_03841_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08182_ (.A1(_03840_),
    .A2(_03841_),
    .ZN(_00922_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08183_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[9] ),
    .A2(_03835_),
    .ZN(_03842_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08184_ (.A1(\u_arbiter.i_wb_cpu_rdt[9] ),
    .A2(_03822_),
    .B1(_03833_),
    .B2(\u_arbiter.i_wb_cpu_dbus_dat[10] ),
    .ZN(_03843_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08185_ (.A1(_03842_),
    .A2(_03843_),
    .ZN(_00923_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08186_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[10] ),
    .A2(_03835_),
    .ZN(_03844_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08187_ (.A1(\u_arbiter.i_wb_cpu_rdt[10] ),
    .A2(_03822_),
    .B1(_03833_),
    .B2(\u_arbiter.i_wb_cpu_dbus_dat[11] ),
    .ZN(_03845_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08188_ (.A1(_03844_),
    .A2(_03845_),
    .ZN(_00924_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08189_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[11] ),
    .A2(_03835_),
    .ZN(_03846_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08190_ (.A1(\u_arbiter.i_wb_cpu_rdt[11] ),
    .A2(_03822_),
    .B1(_03833_),
    .B2(\u_arbiter.i_wb_cpu_dbus_dat[12] ),
    .ZN(_03847_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08191_ (.A1(_03846_),
    .A2(_03847_),
    .ZN(_00925_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08192_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[12] ),
    .A2(_03835_),
    .ZN(_03848_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08193_ (.A1(\u_arbiter.i_wb_cpu_rdt[12] ),
    .A2(_03822_),
    .B1(_03833_),
    .B2(\u_arbiter.i_wb_cpu_dbus_dat[13] ),
    .ZN(_03849_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08194_ (.A1(_03848_),
    .A2(_03849_),
    .ZN(_00926_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08195_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[13] ),
    .A2(_03835_),
    .ZN(_03850_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08196_ (.A1(\u_arbiter.i_wb_cpu_rdt[13] ),
    .A2(_03822_),
    .B1(_03833_),
    .B2(\u_arbiter.i_wb_cpu_dbus_dat[14] ),
    .ZN(_03851_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08197_ (.A1(_03850_),
    .A2(_03851_),
    .ZN(_00927_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08198_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[14] ),
    .A2(_03835_),
    .ZN(_03852_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08199_ (.A1(\u_arbiter.i_wb_cpu_rdt[14] ),
    .A2(_03822_),
    .B1(_03833_),
    .B2(\u_arbiter.i_wb_cpu_dbus_dat[15] ),
    .ZN(_03853_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08200_ (.A1(_03852_),
    .A2(_03853_),
    .ZN(_00928_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08201_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[15] ),
    .A2(_03835_),
    .ZN(_03854_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08202_ (.A1(\u_arbiter.i_wb_cpu_rdt[15] ),
    .A2(_03822_),
    .B1(_03833_),
    .B2(\u_arbiter.i_wb_cpu_dbus_dat[16] ),
    .ZN(_03855_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08203_ (.A1(_03854_),
    .A2(_03855_),
    .ZN(_00929_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08204_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[16] ),
    .A2(_03835_),
    .ZN(_03856_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08205_ (.A1(\u_arbiter.i_wb_cpu_rdt[16] ),
    .A2(_03822_),
    .B1(_03833_),
    .B2(\u_arbiter.i_wb_cpu_dbus_dat[17] ),
    .ZN(_03857_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08206_ (.A1(_03856_),
    .A2(_03857_),
    .ZN(_00930_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08207_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[17] ),
    .A2(_03835_),
    .ZN(_03858_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08208_ (.A1(\u_arbiter.i_wb_cpu_rdt[17] ),
    .A2(_03822_),
    .B1(_03833_),
    .B2(\u_arbiter.i_wb_cpu_dbus_dat[18] ),
    .ZN(_03859_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08209_ (.A1(_03858_),
    .A2(_03859_),
    .ZN(_00931_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08210_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[18] ),
    .A2(_03835_),
    .ZN(_03860_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08211_ (.A1(\u_arbiter.i_wb_cpu_rdt[18] ),
    .A2(_03822_),
    .B1(_03833_),
    .B2(\u_arbiter.i_wb_cpu_dbus_dat[19] ),
    .ZN(_03861_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08212_ (.A1(_03860_),
    .A2(_03861_),
    .ZN(_00932_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08213_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[19] ),
    .A2(_03808_),
    .ZN(_03862_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08214_ (.A1(\u_arbiter.i_wb_cpu_rdt[19] ),
    .A2(_03807_),
    .B1(_03829_),
    .B2(\u_arbiter.i_wb_cpu_dbus_dat[20] ),
    .ZN(_03863_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08215_ (.A1(_03862_),
    .A2(_03863_),
    .ZN(_00933_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08216_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[20] ),
    .A2(_03808_),
    .ZN(_03864_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08217_ (.A1(\u_arbiter.i_wb_cpu_rdt[20] ),
    .A2(_03807_),
    .B1(_03829_),
    .B2(\u_arbiter.i_wb_cpu_dbus_dat[21] ),
    .ZN(_03865_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08218_ (.A1(_03864_),
    .A2(_03865_),
    .ZN(_00934_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08219_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[21] ),
    .A2(_03808_),
    .ZN(_03866_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08220_ (.A1(\u_arbiter.i_wb_cpu_rdt[21] ),
    .A2(_03807_),
    .B1(_03829_),
    .B2(\u_arbiter.i_wb_cpu_dbus_dat[22] ),
    .ZN(_03867_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08221_ (.A1(_03866_),
    .A2(_03867_),
    .ZN(_00935_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08222_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[22] ),
    .A2(_03808_),
    .ZN(_03868_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08223_ (.A1(\u_arbiter.i_wb_cpu_rdt[22] ),
    .A2(_03807_),
    .B1(_03829_),
    .B2(\u_arbiter.i_wb_cpu_dbus_dat[23] ),
    .ZN(_03869_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08224_ (.A1(_03868_),
    .A2(_03869_),
    .ZN(_00936_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08225_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[23] ),
    .A2(_03808_),
    .ZN(_03870_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08226_ (.A1(\u_arbiter.i_wb_cpu_rdt[23] ),
    .A2(_03807_),
    .B1(_03829_),
    .B2(\u_arbiter.i_wb_cpu_dbus_dat[24] ),
    .ZN(_03871_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08227_ (.A1(_03870_),
    .A2(_03871_),
    .ZN(_00937_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08228_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[25] ),
    .A2(_03833_),
    .ZN(_03872_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08229_ (.A1(\u_arbiter.i_wb_cpu_rdt[24] ),
    .A2(_03807_),
    .B1(_03808_),
    .B2(\u_arbiter.i_wb_cpu_dbus_dat[24] ),
    .ZN(_03873_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08230_ (.A1(_03872_),
    .A2(_03873_),
    .ZN(_00938_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08231_ (.A1(_02924_),
    .A2(_03802_),
    .ZN(_03874_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08232_ (.A1(\u_arbiter.i_wb_cpu_rdt[25] ),
    .A2(_03807_),
    .B1(_03808_),
    .B2(\u_arbiter.i_wb_cpu_dbus_dat[25] ),
    .ZN(_03875_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08233_ (.A1(_02445_),
    .A2(_03874_),
    .B(_03875_),
    .ZN(_00939_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _08234_ (.A1(\u_arbiter.i_wb_cpu_rdt[26] ),
    .A2(_02924_),
    .B1(_03874_),
    .B2(\u_arbiter.i_wb_cpu_dbus_dat[27] ),
    .ZN(_03876_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08235_ (.A1(_02445_),
    .A2(_03835_),
    .B(_03876_),
    .ZN(_00940_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08236_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[27] ),
    .A2(_03808_),
    .ZN(_03877_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08237_ (.A1(\u_arbiter.i_wb_cpu_rdt[27] ),
    .A2(_03807_),
    .B1(_03829_),
    .B2(\u_arbiter.i_wb_cpu_dbus_dat[28] ),
    .ZN(_03878_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08238_ (.A1(_03877_),
    .A2(_03878_),
    .ZN(_00941_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08239_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[28] ),
    .A2(_03808_),
    .ZN(_03879_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08240_ (.A1(\u_arbiter.i_wb_cpu_rdt[28] ),
    .A2(_03807_),
    .B1(_03829_),
    .B2(\u_arbiter.i_wb_cpu_dbus_dat[29] ),
    .ZN(_03880_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08241_ (.A1(_03879_),
    .A2(_03880_),
    .ZN(_00942_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08242_ (.A1(\u_arbiter.i_wb_cpu_rdt[29] ),
    .A2(_03807_),
    .B1(_03808_),
    .B2(\u_arbiter.i_wb_cpu_dbus_dat[29] ),
    .ZN(_03881_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08243_ (.A1(_02450_),
    .A2(_03874_),
    .B(_03881_),
    .ZN(_00943_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08244_ (.A1(\u_arbiter.i_wb_cpu_rdt[30] ),
    .A2(_02924_),
    .ZN(_03882_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _08245_ (.A1(_02450_),
    .A2(_03835_),
    .B1(_03833_),
    .B2(_02452_),
    .C(_03882_),
    .ZN(_00944_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _08246_ (.A1(\u_arbiter.i_wb_cpu_rdt[31] ),
    .A2(_02924_),
    .B1(_03874_),
    .B2(_02277_),
    .ZN(_03883_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08247_ (.A1(_02452_),
    .A2(_03835_),
    .B(_03883_),
    .ZN(_00945_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08248_ (.A1(_02695_),
    .A2(_02965_),
    .ZN(_03884_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08249_ (.I(_03884_),
    .Z(_03885_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08250_ (.A1(\u_cpu.rf_ram.memory[113][0] ),
    .A2(_03885_),
    .ZN(_03886_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08251_ (.A1(_03691_),
    .A2(_03885_),
    .B(_03886_),
    .ZN(_00946_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08252_ (.A1(\u_cpu.rf_ram.memory[113][1] ),
    .A2(_03885_),
    .ZN(_03887_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08253_ (.A1(_03695_),
    .A2(_03885_),
    .B(_03887_),
    .ZN(_00947_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08254_ (.A1(\u_cpu.rf_ram.memory[113][2] ),
    .A2(_03885_),
    .ZN(_03888_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08255_ (.A1(_03697_),
    .A2(_03885_),
    .B(_03888_),
    .ZN(_00948_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08256_ (.A1(\u_cpu.rf_ram.memory[113][3] ),
    .A2(_03885_),
    .ZN(_03889_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08257_ (.A1(_03699_),
    .A2(_03885_),
    .B(_03889_),
    .ZN(_00949_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08258_ (.A1(\u_cpu.rf_ram.memory[113][4] ),
    .A2(_03885_),
    .ZN(_03890_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08259_ (.A1(_03701_),
    .A2(_03885_),
    .B(_03890_),
    .ZN(_00950_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08260_ (.A1(\u_cpu.rf_ram.memory[113][5] ),
    .A2(_03885_),
    .ZN(_03891_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08261_ (.A1(_03703_),
    .A2(_03885_),
    .B(_03891_),
    .ZN(_00951_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08262_ (.A1(\u_cpu.rf_ram.memory[113][6] ),
    .A2(_03885_),
    .ZN(_03892_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08263_ (.A1(_03705_),
    .A2(_03885_),
    .B(_03892_),
    .ZN(_00952_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08264_ (.A1(\u_cpu.rf_ram.memory[113][7] ),
    .A2(_03885_),
    .ZN(_03893_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08265_ (.A1(_03707_),
    .A2(_03885_),
    .B(_03893_),
    .ZN(_00953_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08266_ (.A1(_02909_),
    .A2(\u_arbiter.i_wb_cpu_ibus_adr[1] ),
    .ZN(_03894_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08267_ (.A1(\u_arbiter.i_wb_cpu_ack ),
    .A2(_02461_),
    .A3(_03894_),
    .ZN(_03895_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08268_ (.I(_03895_),
    .Z(_03896_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08269_ (.I(_03896_),
    .Z(_03897_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08270_ (.A1(_02465_),
    .A2(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[2] ),
    .ZN(_03898_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08271_ (.A1(_02465_),
    .A2(_02414_),
    .B(_03898_),
    .ZN(_03899_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08272_ (.I0(\u_arbiter.i_wb_cpu_rdt[0] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[0] ),
    .S(_02465_),
    .Z(_03900_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08273_ (.I(_03900_),
    .Z(_03901_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08274_ (.A1(_02465_),
    .A2(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[1] ),
    .ZN(_03902_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08275_ (.A1(_02465_),
    .A2(_02411_),
    .B(_03902_),
    .ZN(_03903_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08276_ (.A1(_03901_),
    .A2(_03903_),
    .ZN(_03904_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08277_ (.I0(\u_arbiter.i_wb_cpu_rdt[14] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[14] ),
    .S(_02465_),
    .Z(_03905_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08278_ (.I(_03905_),
    .Z(_03906_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08279_ (.A1(_02465_),
    .A2(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[15] ),
    .Z(_03907_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08280_ (.A1(_02909_),
    .A2(\u_arbiter.i_wb_cpu_rdt[15] ),
    .B(_03907_),
    .ZN(_03908_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08281_ (.A1(_03906_),
    .A2(_03908_),
    .ZN(_03909_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08282_ (.A1(_03901_),
    .A2(_03903_),
    .ZN(_03910_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08283_ (.A1(_03909_),
    .A2(_03910_),
    .ZN(_03911_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08284_ (.A1(_03904_),
    .A2(_03911_),
    .ZN(_03912_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08285_ (.A1(_02465_),
    .A2(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[0] ),
    .Z(_03913_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08286_ (.A1(_02909_),
    .A2(\u_arbiter.i_wb_cpu_rdt[0] ),
    .B(_03913_),
    .ZN(_03914_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08287_ (.A1(_03914_),
    .A2(_03903_),
    .ZN(_03915_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08288_ (.A1(_02465_),
    .A2(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[13] ),
    .Z(_03916_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08289_ (.A1(_02909_),
    .A2(\u_arbiter.i_wb_cpu_rdt[13] ),
    .B(_03916_),
    .ZN(_03917_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08290_ (.A1(_03906_),
    .A2(_03917_),
    .ZN(_03918_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08291_ (.A1(_03906_),
    .A2(_03908_),
    .ZN(_03919_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08292_ (.I(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[11] ),
    .ZN(_03920_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08293_ (.A1(_02464_),
    .A2(\u_arbiter.i_wb_cpu_rdt[11] ),
    .ZN(_03921_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08294_ (.A1(_02464_),
    .A2(_03920_),
    .B(_03921_),
    .ZN(_03922_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08295_ (.I0(\u_arbiter.i_wb_cpu_rdt[10] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[10] ),
    .S(_02464_),
    .Z(_03923_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08296_ (.I0(\u_arbiter.i_wb_cpu_rdt[9] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[9] ),
    .S(_02464_),
    .Z(_03924_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08297_ (.I0(\u_arbiter.i_wb_cpu_rdt[7] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[7] ),
    .S(_02464_),
    .Z(_03925_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _08298_ (.A1(_03922_),
    .A2(_03923_),
    .A3(_03924_),
    .A4(_03925_),
    .Z(_03926_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08299_ (.A1(_02464_),
    .A2(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[8] ),
    .Z(_03927_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08300_ (.A1(_02909_),
    .A2(\u_arbiter.i_wb_cpu_rdt[8] ),
    .B(_03927_),
    .ZN(_03928_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08301_ (.A1(_03926_),
    .A2(_03928_),
    .ZN(_03929_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _08302_ (.A1(_03917_),
    .A2(_03919_),
    .A3(_03929_),
    .ZN(_03930_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _08303_ (.A1(_03918_),
    .A2(_03930_),
    .Z(_03931_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08304_ (.I0(\u_arbiter.i_wb_cpu_rdt[8] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[8] ),
    .S(_02466_),
    .Z(_03932_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _08305_ (.A1(_03926_),
    .A2(_03932_),
    .Z(_03933_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08306_ (.A1(_02466_),
    .A2(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[12] ),
    .Z(_03934_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08307_ (.A1(_02909_),
    .A2(\u_arbiter.i_wb_cpu_rdt[12] ),
    .B(_03934_),
    .ZN(_03935_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08308_ (.A1(_03933_),
    .A2(_03935_),
    .ZN(_03936_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08309_ (.A1(_02466_),
    .A2(_02411_),
    .ZN(_03937_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08310_ (.A1(_02466_),
    .A2(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[1] ),
    .B(_03937_),
    .ZN(_03938_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08311_ (.A1(_03901_),
    .A2(_03938_),
    .ZN(_03939_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08312_ (.I0(\u_arbiter.i_wb_cpu_rdt[6] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[6] ),
    .S(_02465_),
    .Z(_03940_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08313_ (.I0(\u_arbiter.i_wb_cpu_rdt[5] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[5] ),
    .S(_02465_),
    .Z(_03941_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _08314_ (.A1(_03940_),
    .A2(_03941_),
    .Z(_03942_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08315_ (.A1(_02465_),
    .A2(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[3] ),
    .ZN(_03943_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08316_ (.A1(_02465_),
    .A2(_02416_),
    .B(_03943_),
    .ZN(_03944_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08317_ (.I0(\u_arbiter.i_wb_cpu_rdt[4] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[4] ),
    .S(_02466_),
    .Z(_03945_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _08318_ (.A1(_03942_),
    .A2(_03944_),
    .A3(_03945_),
    .A4(_03899_),
    .ZN(_03946_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08319_ (.I0(\u_arbiter.i_wb_cpu_rdt[15] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[15] ),
    .S(_02465_),
    .Z(_03947_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08320_ (.A1(_03946_),
    .A2(_03947_),
    .ZN(_03948_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08321_ (.A1(_03906_),
    .A2(_03948_),
    .ZN(_03949_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08322_ (.A1(_03939_),
    .A2(_03949_),
    .ZN(_03950_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08323_ (.A1(_03936_),
    .A2(_03950_),
    .ZN(_03951_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _08324_ (.A1(_03899_),
    .A2(_03912_),
    .B1(_03915_),
    .B2(_03931_),
    .C(_03951_),
    .ZN(_03952_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08325_ (.A1(_02265_),
    .A2(_03897_),
    .ZN(_03953_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08326_ (.A1(_03897_),
    .A2(_03952_),
    .B(_03953_),
    .ZN(_00954_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _08327_ (.A1(_03944_),
    .A2(_03912_),
    .B1(_03915_),
    .B2(_03918_),
    .C(_03896_),
    .ZN(_03954_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08328_ (.A1(_02328_),
    .A2(_03897_),
    .B(_03954_),
    .ZN(_00955_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08329_ (.I(_02911_),
    .Z(_03955_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08330_ (.I(_03955_),
    .Z(_03956_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08331_ (.A1(_02466_),
    .A2(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[4] ),
    .Z(_03957_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08332_ (.A1(_02909_),
    .A2(\u_arbiter.i_wb_cpu_rdt[4] ),
    .B(_03957_),
    .ZN(_03958_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08333_ (.A1(_02911_),
    .A2(_03912_),
    .ZN(_03959_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _08334_ (.A1(_03936_),
    .A2(_03938_),
    .A3(_03948_),
    .Z(_03960_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08335_ (.A1(_03914_),
    .A2(_03906_),
    .ZN(_03961_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08336_ (.A1(_03906_),
    .A2(_03947_),
    .ZN(_03962_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08337_ (.A1(_03906_),
    .A2(_03917_),
    .B(_03962_),
    .ZN(_03963_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08338_ (.A1(_03904_),
    .A2(_03911_),
    .Z(_03964_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08339_ (.I(_03964_),
    .Z(_03965_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08340_ (.A1(_02911_),
    .A2(_03965_),
    .ZN(_03966_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08341_ (.A1(_03901_),
    .A2(_03963_),
    .B(_03966_),
    .ZN(_03967_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08342_ (.A1(_03960_),
    .A2(_03961_),
    .A3(_03967_),
    .ZN(_03968_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _08343_ (.A1(_02313_),
    .A2(_03956_),
    .B1(_03958_),
    .B2(_03959_),
    .C(_03968_),
    .ZN(_00956_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08344_ (.A1(_03901_),
    .A2(_03938_),
    .ZN(_03969_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08345_ (.A1(_03909_),
    .A2(_03917_),
    .ZN(_03970_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08346_ (.A1(_03922_),
    .A2(_03923_),
    .ZN(_03971_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08347_ (.I0(\u_arbiter.i_wb_cpu_rdt[13] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[13] ),
    .S(_02466_),
    .Z(_03972_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08348_ (.A1(_02465_),
    .A2(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[14] ),
    .Z(_03973_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08349_ (.A1(_02909_),
    .A2(\u_arbiter.i_wb_cpu_rdt[14] ),
    .B(_03973_),
    .ZN(_03974_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08350_ (.A1(_03974_),
    .A2(_03947_),
    .ZN(_03975_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08351_ (.A1(_03926_),
    .A2(_03928_),
    .B(_03972_),
    .C(_03975_),
    .ZN(_03976_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08352_ (.I(_03963_),
    .ZN(_03977_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08353_ (.A1(_03970_),
    .A2(_03971_),
    .B(_03976_),
    .C(_03977_),
    .ZN(_03978_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08354_ (.A1(_02466_),
    .A2(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[5] ),
    .Z(_03979_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08355_ (.A1(_02909_),
    .A2(\u_arbiter.i_wb_cpu_rdt[5] ),
    .B(_03979_),
    .ZN(_03980_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _08356_ (.A1(_03914_),
    .A2(_03908_),
    .B1(_03912_),
    .B2(_03980_),
    .C(_03896_),
    .ZN(_03981_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08357_ (.A1(_03969_),
    .A2(_03978_),
    .B(_03981_),
    .ZN(_03982_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08358_ (.A1(_02400_),
    .A2(_03956_),
    .B(_03982_),
    .ZN(_00957_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _08359_ (.A1(_02305_),
    .A2(_03956_),
    .B1(_03940_),
    .B2(_03959_),
    .ZN(_03983_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08360_ (.A1(_03950_),
    .A2(_03967_),
    .B(_03983_),
    .ZN(_00958_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08361_ (.A1(_03915_),
    .A2(_03918_),
    .B(_03912_),
    .ZN(_03984_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08362_ (.A1(_03974_),
    .A2(_03908_),
    .ZN(_03985_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08363_ (.A1(_03914_),
    .A2(_03903_),
    .ZN(_03986_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08364_ (.A1(_03940_),
    .A2(_03941_),
    .B(_03971_),
    .ZN(_03987_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08365_ (.A1(_03974_),
    .A2(_03908_),
    .ZN(_03988_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08366_ (.A1(_03899_),
    .A2(_03930_),
    .B1(_03988_),
    .B2(_03972_),
    .ZN(_03989_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08367_ (.A1(_03970_),
    .A2(_03987_),
    .B(_03989_),
    .ZN(_03990_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08368_ (.A1(_03915_),
    .A2(_03990_),
    .ZN(_03991_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _08369_ (.A1(_03935_),
    .A2(_03984_),
    .B1(_03985_),
    .B2(_03986_),
    .C(_03991_),
    .ZN(_03992_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08370_ (.A1(_03956_),
    .A2(_03992_),
    .ZN(_03993_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08371_ (.A1(_02286_),
    .A2(_03956_),
    .B(_03993_),
    .ZN(_00959_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08372_ (.A1(_03965_),
    .A2(_03961_),
    .ZN(_03994_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08373_ (.A1(_02466_),
    .A2(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[10] ),
    .Z(_03995_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08374_ (.A1(_02909_),
    .A2(\u_arbiter.i_wb_cpu_rdt[10] ),
    .B(_03995_),
    .ZN(_03996_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08375_ (.A1(_03974_),
    .A2(_03947_),
    .ZN(_03997_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08376_ (.A1(_03997_),
    .A2(_03972_),
    .ZN(_03998_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08377_ (.A1(_03996_),
    .A2(_03940_),
    .B(_03998_),
    .C(_03922_),
    .ZN(_03999_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08378_ (.I0(\u_arbiter.i_wb_cpu_rdt[12] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[12] ),
    .S(_02466_),
    .Z(_04000_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08379_ (.A1(_04000_),
    .A2(_03918_),
    .B1(_03930_),
    .B2(_03944_),
    .ZN(_04001_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08380_ (.A1(_03999_),
    .A2(_04001_),
    .B(_03969_),
    .ZN(_04002_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _08381_ (.A1(_03965_),
    .A2(_03972_),
    .B1(_03994_),
    .B2(_04002_),
    .C(_03955_),
    .ZN(_04003_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08382_ (.A1(_02285_),
    .A2(_03956_),
    .B(_04003_),
    .ZN(_00960_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08383_ (.A1(_03942_),
    .A2(_03971_),
    .ZN(_04004_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08384_ (.A1(_03970_),
    .A2(_04004_),
    .ZN(_04005_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _08385_ (.A1(_04000_),
    .A2(_03918_),
    .B1(_03930_),
    .B2(_03945_),
    .C(_04005_),
    .ZN(_04006_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _08386_ (.A1(_03974_),
    .A2(_03904_),
    .B1(_03969_),
    .B2(_04006_),
    .ZN(_04007_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08387_ (.A1(_03956_),
    .A2(_04007_),
    .ZN(_04008_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08388_ (.A1(_02309_),
    .A2(_03956_),
    .B(_04008_),
    .ZN(_00961_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08389_ (.A1(_03895_),
    .A2(_03965_),
    .ZN(_04009_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08390_ (.I0(\u_arbiter.i_wb_cpu_rdt[20] ),
    .I1(\u_arbiter.i_wb_cpu_rdt[4] ),
    .S(_02467_),
    .Z(_04010_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _08391_ (.A1(_03936_),
    .A2(_03949_),
    .B1(_03919_),
    .B2(_03899_),
    .C(_03938_),
    .ZN(_04011_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08392_ (.A1(_03899_),
    .A2(_03917_),
    .A3(_03962_),
    .ZN(_04012_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08393_ (.A1(_04000_),
    .A2(_03931_),
    .ZN(_04013_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08394_ (.A1(_03901_),
    .A2(_04012_),
    .A3(_04013_),
    .ZN(_04014_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08395_ (.A1(_03899_),
    .A2(_03988_),
    .ZN(_04015_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08396_ (.A1(_03910_),
    .A2(_04015_),
    .ZN(_04016_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _08397_ (.A1(_02911_),
    .A2(_03904_),
    .A3(_04014_),
    .A4(_04016_),
    .ZN(_04017_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08398_ (.A1(_04011_),
    .A2(_04017_),
    .ZN(_04018_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08399_ (.A1(_04009_),
    .A2(_04010_),
    .B(_04018_),
    .ZN(_04019_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08400_ (.A1(_02325_),
    .A2(_03956_),
    .B(_04019_),
    .ZN(_00962_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08401_ (.I0(\u_arbiter.i_wb_cpu_rdt[21] ),
    .I1(\u_arbiter.i_wb_cpu_rdt[5] ),
    .S(_02467_),
    .Z(_04020_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08402_ (.A1(_03944_),
    .A2(_03988_),
    .ZN(_04021_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08403_ (.A1(_04000_),
    .A2(_03930_),
    .ZN(_04022_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08404_ (.A1(_03901_),
    .A2(_04022_),
    .ZN(_04023_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08405_ (.A1(_03947_),
    .A2(_03972_),
    .ZN(_04024_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08406_ (.A1(_03974_),
    .A2(_04024_),
    .B(_03938_),
    .ZN(_04025_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08407_ (.A1(_03901_),
    .A2(_03975_),
    .B(_04025_),
    .ZN(_04026_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08408_ (.A1(_03938_),
    .A2(_04023_),
    .B1(_04026_),
    .B2(_03944_),
    .ZN(_04027_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08409_ (.A1(_03910_),
    .A2(_04021_),
    .B(_04027_),
    .ZN(_04028_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08410_ (.A1(_04009_),
    .A2(_04020_),
    .B1(_04028_),
    .B2(_03955_),
    .ZN(_04029_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08411_ (.A1(_01448_),
    .A2(_03956_),
    .B(_04029_),
    .ZN(_00963_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08412_ (.I0(\u_arbiter.i_wb_cpu_rdt[22] ),
    .I1(\u_arbiter.i_wb_cpu_rdt[6] ),
    .S(_02466_),
    .Z(_04030_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08413_ (.A1(_03914_),
    .A2(_03938_),
    .ZN(_04031_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _08414_ (.A1(_03940_),
    .A2(_03908_),
    .B1(_03909_),
    .B2(_04030_),
    .C1(_03988_),
    .C2(_03945_),
    .ZN(_04032_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08415_ (.A1(_03935_),
    .A2(_03976_),
    .ZN(_04033_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _08416_ (.A1(_03974_),
    .A2(_04033_),
    .A3(_04024_),
    .B(_03915_),
    .ZN(_04034_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08417_ (.A1(_03986_),
    .A2(_04034_),
    .ZN(_04035_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08418_ (.A1(_03969_),
    .A2(_04022_),
    .B(_03958_),
    .ZN(_04036_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08419_ (.A1(_04035_),
    .A2(_04036_),
    .ZN(_04037_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08420_ (.A1(_04031_),
    .A2(_04032_),
    .B(_04037_),
    .C(_03965_),
    .ZN(_04038_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08421_ (.A1(_03965_),
    .A2(_04030_),
    .B(_04038_),
    .C(_03955_),
    .ZN(_04039_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08422_ (.A1(_02290_),
    .A2(_03956_),
    .B(_04039_),
    .ZN(_00964_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08423_ (.A1(_02619_),
    .A2(_02965_),
    .ZN(_04040_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08424_ (.I(_04040_),
    .Z(_04041_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08425_ (.A1(\u_cpu.rf_ram.memory[114][0] ),
    .A2(_04041_),
    .ZN(_04042_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08426_ (.A1(_03691_),
    .A2(_04041_),
    .B(_04042_),
    .ZN(_00965_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08427_ (.A1(\u_cpu.rf_ram.memory[114][1] ),
    .A2(_04041_),
    .ZN(_04043_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08428_ (.A1(_03695_),
    .A2(_04041_),
    .B(_04043_),
    .ZN(_00966_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08429_ (.A1(\u_cpu.rf_ram.memory[114][2] ),
    .A2(_04041_),
    .ZN(_04044_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08430_ (.A1(_03697_),
    .A2(_04041_),
    .B(_04044_),
    .ZN(_00967_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08431_ (.A1(\u_cpu.rf_ram.memory[114][3] ),
    .A2(_04041_),
    .ZN(_04045_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08432_ (.A1(_03699_),
    .A2(_04041_),
    .B(_04045_),
    .ZN(_00968_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08433_ (.A1(\u_cpu.rf_ram.memory[114][4] ),
    .A2(_04041_),
    .ZN(_04046_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08434_ (.A1(_03701_),
    .A2(_04041_),
    .B(_04046_),
    .ZN(_00969_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08435_ (.A1(\u_cpu.rf_ram.memory[114][5] ),
    .A2(_04041_),
    .ZN(_04047_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08436_ (.A1(_03703_),
    .A2(_04041_),
    .B(_04047_),
    .ZN(_00970_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08437_ (.A1(\u_cpu.rf_ram.memory[114][6] ),
    .A2(_04041_),
    .ZN(_04048_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08438_ (.A1(_03705_),
    .A2(_04041_),
    .B(_04048_),
    .ZN(_00971_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08439_ (.A1(\u_cpu.rf_ram.memory[114][7] ),
    .A2(_04041_),
    .ZN(_04049_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08440_ (.A1(_03707_),
    .A2(_04041_),
    .B(_04049_),
    .ZN(_00972_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08441_ (.I0(\u_arbiter.i_wb_cpu_rdt[26] ),
    .I1(\u_arbiter.i_wb_cpu_rdt[10] ),
    .S(_02466_),
    .Z(_04050_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08442_ (.A1(_03906_),
    .A2(_03947_),
    .ZN(_04051_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08443_ (.A1(_03917_),
    .A2(_04051_),
    .ZN(_04052_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08444_ (.A1(_04000_),
    .A2(_04052_),
    .B(_03915_),
    .ZN(_04053_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08445_ (.A1(_03935_),
    .A2(_03974_),
    .ZN(_04054_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _08446_ (.A1(_03922_),
    .A2(_03996_),
    .A3(_04000_),
    .A4(_03998_),
    .Z(_04055_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08447_ (.A1(_04024_),
    .A2(_04054_),
    .B(_04055_),
    .ZN(_04056_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08448_ (.A1(_04052_),
    .A2(_04056_),
    .ZN(_04057_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08449_ (.A1(_04000_),
    .A2(_03929_),
    .B(_03975_),
    .C(_03972_),
    .ZN(_04058_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08450_ (.A1(_03980_),
    .A2(_03929_),
    .B(_04058_),
    .ZN(_04059_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08451_ (.A1(_03925_),
    .A2(_03918_),
    .B1(_03988_),
    .B2(_03941_),
    .ZN(_04060_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08452_ (.I(_04060_),
    .ZN(_04061_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _08453_ (.A1(_04057_),
    .A2(_04059_),
    .A3(_04061_),
    .ZN(_04062_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _08454_ (.A1(_03899_),
    .A2(_03975_),
    .B1(_03988_),
    .B2(_03925_),
    .C(_03938_),
    .ZN(_04063_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _08455_ (.A1(_04053_),
    .A2(_04062_),
    .B1(_04063_),
    .B2(_03901_),
    .ZN(_04064_));
 gf180mcu_fd_sc_mcu7t5v0__oai222_1 _08456_ (.A1(_03974_),
    .A2(_03941_),
    .B1(_03997_),
    .B2(_04050_),
    .C1(_03985_),
    .C2(_03925_),
    .ZN(_04065_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08457_ (.A1(_03910_),
    .A2(_04065_),
    .B(_03966_),
    .ZN(_04066_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08458_ (.A1(_04009_),
    .A2(_04050_),
    .B1(_04064_),
    .B2(_04066_),
    .ZN(_04067_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08459_ (.A1(_01454_),
    .A2(_03956_),
    .B(_04067_),
    .ZN(_00973_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _08460_ (.A1(_02265_),
    .A2(_02400_),
    .A3(_01446_),
    .B(_02259_),
    .ZN(_04068_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08461_ (.A1(_03896_),
    .A2(_04068_),
    .Z(_04069_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08462_ (.A1(_03955_),
    .A2(_04068_),
    .ZN(_04070_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08463_ (.A1(\u_cpu.cpu.immdec.imm24_20[0] ),
    .A2(_04069_),
    .B1(_04070_),
    .B2(\u_cpu.cpu.immdec.imm24_20[1] ),
    .ZN(_04071_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08464_ (.A1(_04019_),
    .A2(_04071_),
    .ZN(_00974_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08465_ (.A1(\u_cpu.cpu.immdec.imm24_20[1] ),
    .A2(_04069_),
    .B1(_04070_),
    .B2(\u_cpu.cpu.immdec.imm24_20[2] ),
    .ZN(_04072_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08466_ (.A1(_04029_),
    .A2(_04072_),
    .ZN(_00975_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08467_ (.I(\u_cpu.cpu.immdec.imm24_20[2] ),
    .ZN(_04073_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08468_ (.A1(\u_cpu.cpu.immdec.imm24_20[3] ),
    .A2(_04068_),
    .B(_03896_),
    .ZN(_04074_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08469_ (.A1(_04073_),
    .A2(_04069_),
    .B1(_04074_),
    .B2(_04039_),
    .ZN(_00976_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08470_ (.I0(\u_arbiter.i_wb_cpu_rdt[23] ),
    .I1(\u_arbiter.i_wb_cpu_rdt[7] ),
    .S(_02466_),
    .Z(_04075_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08471_ (.A1(_03970_),
    .A2(_03971_),
    .B(_04022_),
    .ZN(_04076_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08472_ (.I(_04034_),
    .ZN(_04077_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08473_ (.A1(_03941_),
    .A2(_04035_),
    .B1(_04076_),
    .B2(_04077_),
    .ZN(_04078_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08474_ (.A1(_03996_),
    .A2(_03908_),
    .ZN(_04079_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08475_ (.A1(_03906_),
    .A2(_04079_),
    .ZN(_04080_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _08476_ (.A1(_03941_),
    .A2(_04051_),
    .B1(_04075_),
    .B2(_03947_),
    .C(_04031_),
    .ZN(_04081_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _08477_ (.A1(_04031_),
    .A2(_04078_),
    .B1(_04080_),
    .B2(_04081_),
    .C(_03912_),
    .ZN(_04082_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08478_ (.A1(_03912_),
    .A2(_04075_),
    .B(_04082_),
    .C(_03896_),
    .ZN(_04083_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08479_ (.A1(\u_cpu.cpu.immdec.imm24_20[4] ),
    .A2(_03955_),
    .ZN(_04084_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08480_ (.A1(\u_cpu.cpu.immdec.imm24_20[3] ),
    .A2(_04069_),
    .ZN(_04085_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _08481_ (.A1(_04069_),
    .A2(_04083_),
    .A3(_04084_),
    .B(_04085_),
    .ZN(_00977_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08482_ (.I(_03978_),
    .ZN(_04086_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _08483_ (.A1(_03922_),
    .A2(_03918_),
    .B1(_04086_),
    .B2(_03940_),
    .C(_04023_),
    .ZN(_04087_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08484_ (.I0(\u_arbiter.i_wb_cpu_rdt[24] ),
    .I1(\u_arbiter.i_wb_cpu_rdt[8] ),
    .S(_02467_),
    .Z(_04088_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _08485_ (.A1(_03922_),
    .A2(_03908_),
    .B1(_03909_),
    .B2(_04088_),
    .C(_04031_),
    .ZN(_04089_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08486_ (.A1(_03914_),
    .A2(_03940_),
    .B(_03938_),
    .ZN(_04090_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _08487_ (.A1(_03966_),
    .A2(_04087_),
    .A3(_04089_),
    .A4(_04090_),
    .Z(_04091_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _08488_ (.A1(\u_cpu.cpu.immdec.imm24_20[4] ),
    .A2(_04069_),
    .B1(_04070_),
    .B2(\u_cpu.cpu.immdec.imm30_25[0] ),
    .C1(_04088_),
    .C2(_04009_),
    .ZN(_04092_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08489_ (.A1(_04091_),
    .A2(_04092_),
    .ZN(_00978_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _08490_ (.A1(_03926_),
    .A2(_03928_),
    .A3(_03917_),
    .ZN(_04093_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08491_ (.A1(_03963_),
    .A2(_04093_),
    .B(_03899_),
    .ZN(_04094_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08492_ (.A1(_04000_),
    .A2(_04024_),
    .B(_04055_),
    .C(_04033_),
    .ZN(_04095_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08493_ (.A1(_03901_),
    .A2(_04094_),
    .A3(_04095_),
    .ZN(_04096_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08494_ (.A1(_03935_),
    .A2(_03914_),
    .B1(_03903_),
    .B2(_03961_),
    .ZN(_04097_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08495_ (.A1(_04096_),
    .A2(_04097_),
    .B(_03966_),
    .ZN(_04098_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08496_ (.I0(\u_arbiter.i_wb_cpu_rdt[25] ),
    .I1(\u_arbiter.i_wb_cpu_rdt[9] ),
    .S(_02467_),
    .Z(_04099_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _08497_ (.A1(_01444_),
    .A2(_02305_),
    .A3(\u_arbiter.i_wb_cpu_dbus_we ),
    .ZN(_04100_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08498_ (.A1(_02265_),
    .A2(_04100_),
    .B(_02392_),
    .ZN(_04101_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _08499_ (.A1(_03955_),
    .A2(_04101_),
    .Z(_04102_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _08500_ (.A1(\u_cpu.cpu.immdec.imm30_25[1] ),
    .A2(_03956_),
    .B1(_03959_),
    .B2(_04099_),
    .C(_04102_),
    .ZN(_04103_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08501_ (.A1(_03955_),
    .A2(_04101_),
    .ZN(_04104_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08502_ (.A1(\u_cpu.cpu.immdec.imm30_25[0] ),
    .A2(_04104_),
    .ZN(_04105_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08503_ (.A1(_04098_),
    .A2(_04103_),
    .B(_04105_),
    .ZN(_00979_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08504_ (.A1(_03896_),
    .A2(_04101_),
    .Z(_04106_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08505_ (.A1(\u_cpu.cpu.immdec.imm30_25[1] ),
    .A2(_04104_),
    .B1(_04106_),
    .B2(\u_cpu.cpu.immdec.imm30_25[2] ),
    .ZN(_04107_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08506_ (.A1(_04067_),
    .A2(_04107_),
    .ZN(_00980_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08507_ (.A1(_03944_),
    .A2(_03975_),
    .A3(_04093_),
    .ZN(_04108_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08508_ (.A1(_03940_),
    .A2(_03963_),
    .ZN(_04109_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _08509_ (.A1(_03901_),
    .A2(_04095_),
    .A3(_04108_),
    .A4(_04109_),
    .ZN(_04110_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08510_ (.A1(_03932_),
    .A2(_03988_),
    .ZN(_04111_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08511_ (.A1(_03944_),
    .A2(_03975_),
    .B(_03938_),
    .ZN(_04112_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08512_ (.I0(\u_arbiter.i_wb_cpu_rdt[27] ),
    .I1(\u_arbiter.i_wb_cpu_rdt[11] ),
    .S(_02466_),
    .Z(_04113_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08513_ (.A1(_03932_),
    .A2(_04051_),
    .B1(_04113_),
    .B2(_03909_),
    .ZN(_04114_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _08514_ (.A1(_04111_),
    .A2(_04112_),
    .B1(_04114_),
    .B2(_03910_),
    .C(_03966_),
    .ZN(_04115_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08515_ (.A1(_04110_),
    .A2(_04115_),
    .ZN(_04116_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _08516_ (.A1(\u_cpu.cpu.immdec.imm30_25[2] ),
    .A2(_04104_),
    .B1(_04106_),
    .B2(\u_cpu.cpu.immdec.imm30_25[3] ),
    .C1(_04113_),
    .C2(_04009_),
    .ZN(_04117_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08517_ (.A1(_04116_),
    .A2(_04117_),
    .ZN(_00981_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08518_ (.A1(_03924_),
    .A2(_03918_),
    .B1(_03988_),
    .B2(_04000_),
    .ZN(_04118_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08519_ (.A1(_03958_),
    .A2(_03929_),
    .B(_04058_),
    .ZN(_04119_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08520_ (.A1(_04057_),
    .A2(_04119_),
    .ZN(_04120_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08521_ (.A1(_04118_),
    .A2(_04120_),
    .B(_04053_),
    .ZN(_04121_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _08522_ (.A1(_03924_),
    .A2(_03910_),
    .A3(_04051_),
    .Z(_04122_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _08523_ (.A1(_03966_),
    .A2(_04121_),
    .A3(_04122_),
    .ZN(_04123_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08524_ (.A1(_03896_),
    .A2(_04101_),
    .ZN(_04124_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08525_ (.I0(\u_arbiter.i_wb_cpu_rdt[28] ),
    .I1(\u_arbiter.i_wb_cpu_rdt[12] ),
    .S(_02467_),
    .Z(_04125_));
 gf180mcu_fd_sc_mcu7t5v0__oai222_1 _08526_ (.A1(\u_cpu.cpu.immdec.imm30_25[3] ),
    .A2(_04102_),
    .B1(_04124_),
    .B2(\u_cpu.cpu.immdec.imm30_25[4] ),
    .C1(_04125_),
    .C2(_03959_),
    .ZN(_04126_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08527_ (.A1(_04123_),
    .A2(_04126_),
    .ZN(_00982_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08528_ (.A1(_03923_),
    .A2(_03918_),
    .ZN(_04127_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08529_ (.A1(_03935_),
    .A2(_03974_),
    .B(_04052_),
    .ZN(_04128_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08530_ (.A1(_04055_),
    .A2(_04128_),
    .ZN(_04129_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08531_ (.A1(_04127_),
    .A2(_04129_),
    .B(_04053_),
    .ZN(_04130_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08532_ (.I0(\u_arbiter.i_wb_cpu_rdt[29] ),
    .I1(\u_arbiter.i_wb_cpu_rdt[13] ),
    .S(_02467_),
    .Z(_04131_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08533_ (.A1(_03908_),
    .A2(_04131_),
    .B(_04079_),
    .C(_03910_),
    .ZN(_04132_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08534_ (.A1(_03906_),
    .A2(_04132_),
    .ZN(_04133_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _08535_ (.A1(_03966_),
    .A2(_04130_),
    .A3(_04133_),
    .ZN(_04134_));
 gf180mcu_fd_sc_mcu7t5v0__oai222_1 _08536_ (.A1(\u_cpu.cpu.immdec.imm30_25[4] ),
    .A2(_04102_),
    .B1(_04124_),
    .B2(\u_cpu.cpu.immdec.imm30_25[5] ),
    .C1(_04131_),
    .C2(_03959_),
    .ZN(_04135_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08537_ (.A1(_04134_),
    .A2(_04135_),
    .ZN(_00983_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08538_ (.I0(\u_arbiter.i_wb_cpu_rdt[30] ),
    .I1(\u_arbiter.i_wb_cpu_rdt[14] ),
    .S(_02467_),
    .Z(_04136_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08539_ (.A1(_03923_),
    .A2(_03935_),
    .B(_03922_),
    .ZN(_04137_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _08540_ (.A1(_03922_),
    .A2(_03923_),
    .B1(_04004_),
    .B2(_04137_),
    .C(_03998_),
    .ZN(_04138_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08541_ (.A1(_03932_),
    .A2(_03918_),
    .B(_04128_),
    .ZN(_04139_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08542_ (.A1(_04138_),
    .A2(_04139_),
    .B(_04053_),
    .ZN(_04140_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08543_ (.A1(_04009_),
    .A2(_04136_),
    .B1(_04140_),
    .B2(_03955_),
    .ZN(_04141_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08544_ (.A1(\u_cpu.cpu.immdec.imm30_25[5] ),
    .A2(_04104_),
    .ZN(_04142_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08545_ (.I(\u_cpu.cpu.immdec.imm19_12_20[0] ),
    .ZN(_04143_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08546_ (.A1(_01444_),
    .A2(_02265_),
    .B(\u_cpu.cpu.decode.opcode[1] ),
    .ZN(_04144_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08547_ (.A1(_02320_),
    .A2(_04144_),
    .ZN(_04145_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08548_ (.A1(_04143_),
    .A2(_04144_),
    .B(_04145_),
    .C(_02585_),
    .ZN(_04146_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08549_ (.A1(\u_cpu.cpu.immdec.imm7 ),
    .A2(_02585_),
    .B(_04106_),
    .C(_04146_),
    .ZN(_04147_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08550_ (.A1(_04141_),
    .A2(_04142_),
    .A3(_04147_),
    .ZN(_00984_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08551_ (.A1(_03925_),
    .A2(_04052_),
    .ZN(_04148_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08552_ (.A1(_03969_),
    .A2(_04148_),
    .ZN(_04149_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _08553_ (.A1(_03925_),
    .A2(_03974_),
    .Z(_04150_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08554_ (.A1(_03925_),
    .A2(_03998_),
    .B1(_04150_),
    .B2(_03908_),
    .ZN(_04151_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08555_ (.A1(_03935_),
    .A2(_03962_),
    .B(_04151_),
    .ZN(_04152_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08556_ (.A1(_03933_),
    .A2(_04000_),
    .A3(_03949_),
    .ZN(_04153_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08557_ (.A1(_03925_),
    .A2(_03948_),
    .A3(_03962_),
    .ZN(_04154_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08558_ (.A1(_03903_),
    .A2(_04153_),
    .A3(_04154_),
    .ZN(_04155_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08559_ (.A1(_04149_),
    .A2(_04152_),
    .B1(_04155_),
    .B2(_03914_),
    .ZN(_04156_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _08560_ (.A1(_03899_),
    .A2(_03908_),
    .B1(_03909_),
    .B2(_03925_),
    .C(_04031_),
    .ZN(_04157_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08561_ (.A1(_04156_),
    .A2(_04157_),
    .ZN(_04158_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08562_ (.A1(_03896_),
    .A2(_03912_),
    .ZN(_04159_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08563_ (.A1(_03925_),
    .A2(_04009_),
    .B1(_04158_),
    .B2(_04159_),
    .ZN(_04160_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08564_ (.A1(_02392_),
    .A2(_02320_),
    .B(_03896_),
    .ZN(_04161_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08565_ (.A1(\u_cpu.cpu.immdec.imm7 ),
    .A2(_02259_),
    .ZN(_04162_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08566_ (.A1(_04160_),
    .A2(_04161_),
    .B1(_04162_),
    .B2(_03897_),
    .ZN(_00985_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08567_ (.A1(_01444_),
    .A2(_02328_),
    .B(_02269_),
    .C(_02318_),
    .ZN(_04163_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08568_ (.A1(_02259_),
    .A2(_04163_),
    .B(_02911_),
    .ZN(_04164_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08569_ (.I(_04164_),
    .Z(_04165_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08570_ (.A1(\u_cpu.cpu.immdec.imm19_12_20[1] ),
    .A2(_03897_),
    .B(_04165_),
    .ZN(_04166_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08571_ (.A1(_04143_),
    .A2(_04165_),
    .B1(_04166_),
    .B2(_04019_),
    .ZN(_00986_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08572_ (.I(\u_cpu.cpu.immdec.imm19_12_20[1] ),
    .ZN(_04167_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08573_ (.A1(\u_cpu.cpu.immdec.imm19_12_20[2] ),
    .A2(_03897_),
    .B(_04165_),
    .ZN(_04168_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08574_ (.A1(_04167_),
    .A2(_04165_),
    .B1(_04168_),
    .B2(_03993_),
    .ZN(_00987_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08575_ (.I(\u_cpu.cpu.immdec.imm19_12_20[2] ),
    .ZN(_04169_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08576_ (.A1(\u_cpu.cpu.immdec.imm19_12_20[3] ),
    .A2(_03897_),
    .B(_04165_),
    .ZN(_04170_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08577_ (.A1(_04169_),
    .A2(_04165_),
    .B1(_04170_),
    .B2(_04003_),
    .ZN(_00988_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08578_ (.I(\u_cpu.cpu.immdec.imm19_12_20[3] ),
    .ZN(_04171_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08579_ (.A1(\u_cpu.cpu.csr_imm ),
    .A2(_03897_),
    .B(_04164_),
    .ZN(_04172_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08580_ (.A1(_04171_),
    .A2(_04165_),
    .B1(_04172_),
    .B2(_04008_),
    .ZN(_00989_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08581_ (.A1(_04000_),
    .A2(_03918_),
    .ZN(_04173_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08582_ (.A1(_03980_),
    .A2(_03976_),
    .B(_04173_),
    .C(_04052_),
    .ZN(_04174_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08583_ (.A1(_04149_),
    .A2(_04174_),
    .ZN(_04175_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08584_ (.A1(_03910_),
    .A2(_03985_),
    .A3(_04150_),
    .ZN(_04176_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _08585_ (.A1(_04000_),
    .A2(_03946_),
    .A3(_03908_),
    .ZN(_04177_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _08586_ (.A1(_03986_),
    .A2(_03906_),
    .A3(_04177_),
    .ZN(_04178_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08587_ (.A1(_03924_),
    .A2(_04052_),
    .B(_03915_),
    .ZN(_04179_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _08588_ (.A1(_03908_),
    .A2(_03918_),
    .A3(_04179_),
    .ZN(_04180_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08589_ (.A1(_04178_),
    .A2(_04180_),
    .B(_03925_),
    .ZN(_04181_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _08590_ (.A1(_03965_),
    .A2(_04175_),
    .A3(_04176_),
    .A4(_04181_),
    .ZN(_04182_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08591_ (.A1(_03947_),
    .A2(_03904_),
    .B(_04182_),
    .C(_03955_),
    .ZN(_04183_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08592_ (.A1(\u_cpu.cpu.immdec.imm19_12_20[5] ),
    .A2(_03897_),
    .B(_04165_),
    .ZN(_04184_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08593_ (.A1(_01439_),
    .A2(_04165_),
    .B1(_04183_),
    .B2(_04184_),
    .ZN(_00990_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08594_ (.I0(\u_arbiter.i_wb_cpu_rdt[16] ),
    .I1(\u_arbiter.i_wb_cpu_rdt[0] ),
    .S(_02466_),
    .Z(_04185_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08595_ (.A1(_03909_),
    .A2(_04185_),
    .ZN(_04186_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08596_ (.A1(_03932_),
    .A2(_03906_),
    .B(_04031_),
    .C(_04051_),
    .ZN(_04187_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08597_ (.A1(_03972_),
    .A2(_03985_),
    .ZN(_04188_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08598_ (.A1(_03940_),
    .A2(_03929_),
    .B(_03975_),
    .C(_03972_),
    .ZN(_04189_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08599_ (.A1(_03932_),
    .A2(_03998_),
    .ZN(_04190_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _08600_ (.A1(_04173_),
    .A2(_04052_),
    .A3(_04111_),
    .A4(_04190_),
    .Z(_04191_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _08601_ (.A1(_03928_),
    .A2(_04188_),
    .B1(_04189_),
    .B2(_04191_),
    .C(_03969_),
    .ZN(_04192_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _08602_ (.A1(_03928_),
    .A2(_03986_),
    .A3(_04177_),
    .ZN(_04193_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08603_ (.A1(_04031_),
    .A2(_03961_),
    .ZN(_04194_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _08604_ (.A1(_04192_),
    .A2(_04193_),
    .A3(_04194_),
    .ZN(_04195_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08605_ (.A1(_04186_),
    .A2(_04187_),
    .B(_03912_),
    .C(_04195_),
    .ZN(_04196_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08606_ (.A1(_03912_),
    .A2(_04185_),
    .B(_04196_),
    .C(_03896_),
    .ZN(_04197_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08607_ (.A1(\u_cpu.cpu.immdec.imm19_12_20[6] ),
    .A2(_03955_),
    .ZN(_04198_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08608_ (.A1(\u_cpu.cpu.immdec.imm19_12_20[5] ),
    .A2(_04165_),
    .ZN(_04199_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _08609_ (.A1(_04165_),
    .A2(_04197_),
    .A3(_04198_),
    .B(_04199_),
    .ZN(_00991_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08610_ (.A1(\u_cpu.cpu.immdec.imm19_12_20[6] ),
    .A2(_04165_),
    .ZN(_04200_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08611_ (.A1(_02909_),
    .A2(\u_arbiter.i_wb_cpu_rdt[17] ),
    .ZN(_04201_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08612_ (.A1(_02909_),
    .A2(_02411_),
    .B(_04201_),
    .ZN(_04202_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08613_ (.A1(_04013_),
    .A2(_04052_),
    .B(_04179_),
    .ZN(_04203_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08614_ (.A1(_04178_),
    .A2(_04180_),
    .B(_03924_),
    .ZN(_04204_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08615_ (.A1(_04031_),
    .A2(_04204_),
    .ZN(_04205_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08616_ (.A1(_04203_),
    .A2(_04205_),
    .ZN(_04206_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _08617_ (.A1(_03924_),
    .A2(_03906_),
    .B1(_03909_),
    .B2(_04202_),
    .C(_04031_),
    .ZN(_04207_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08618_ (.A1(_04206_),
    .A2(_04207_),
    .B(_04159_),
    .ZN(_04208_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08619_ (.A1(\u_cpu.cpu.immdec.imm19_12_20[7] ),
    .A2(_03955_),
    .ZN(_04209_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08620_ (.A1(_04164_),
    .A2(_04209_),
    .ZN(_04210_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08621_ (.A1(_03959_),
    .A2(_04202_),
    .B(_04208_),
    .C(_04210_),
    .ZN(_04211_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08622_ (.A1(_04200_),
    .A2(_04211_),
    .ZN(_00992_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08623_ (.A1(_03923_),
    .A2(_04178_),
    .B(_03910_),
    .ZN(_04212_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08624_ (.A1(_03918_),
    .A2(_03975_),
    .B(_04013_),
    .ZN(_04213_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08625_ (.A1(_03923_),
    .A2(_04052_),
    .B(_04213_),
    .C(_03915_),
    .ZN(_04214_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08626_ (.A1(_03974_),
    .A2(_03910_),
    .B1(_04212_),
    .B2(_04214_),
    .ZN(_04215_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08627_ (.A1(_02467_),
    .A2(\u_arbiter.i_wb_cpu_rdt[18] ),
    .ZN(_04216_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08628_ (.A1(_02467_),
    .A2(_02414_),
    .B(_03965_),
    .C(_04216_),
    .ZN(_04217_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _08629_ (.A1(_03896_),
    .A2(_04215_),
    .A3(_04217_),
    .ZN(_04218_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08630_ (.A1(\u_cpu.cpu.immdec.imm19_12_20[8] ),
    .A2(_03955_),
    .ZN(_04219_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08631_ (.A1(\u_cpu.cpu.immdec.imm19_12_20[7] ),
    .A2(_04165_),
    .ZN(_04220_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _08632_ (.A1(_04165_),
    .A2(_04218_),
    .A3(_04219_),
    .B(_04220_),
    .ZN(_00993_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08633_ (.A1(_03922_),
    .A2(_04188_),
    .ZN(_04221_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08634_ (.A1(_04013_),
    .A2(_04221_),
    .B(_03969_),
    .ZN(_04222_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08635_ (.A1(_02467_),
    .A2(_02416_),
    .ZN(_04223_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08636_ (.A1(_02467_),
    .A2(\u_arbiter.i_wb_cpu_rdt[19] ),
    .B(_03912_),
    .C(_04223_),
    .ZN(_04224_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08637_ (.A1(_03955_),
    .A2(_04224_),
    .ZN(_04225_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08638_ (.A1(_03922_),
    .A2(_04178_),
    .B(_04222_),
    .C(_04225_),
    .ZN(_04226_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08639_ (.A1(_02305_),
    .A2(_01440_),
    .B(_03896_),
    .ZN(_04227_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08640_ (.A1(_02305_),
    .A2(_02320_),
    .B(_04227_),
    .ZN(_04228_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08641_ (.A1(\u_cpu.cpu.immdec.imm19_12_20[8] ),
    .A2(_04165_),
    .ZN(_04229_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _08642_ (.A1(_04165_),
    .A2(_04226_),
    .A3(_04228_),
    .B(_04229_),
    .ZN(_00994_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08643_ (.I0(\u_arbiter.i_wb_cpu_rdt[31] ),
    .I1(\u_arbiter.i_wb_cpu_rdt[15] ),
    .S(_02467_),
    .Z(_04230_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08644_ (.A1(_04173_),
    .A2(_04129_),
    .B(_04053_),
    .C(_03896_),
    .ZN(_04231_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _08645_ (.A1(\u_cpu.cpu.immdec.imm31 ),
    .A2(_03897_),
    .B1(_04009_),
    .B2(_04230_),
    .C(_04231_),
    .ZN(_04232_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _08646_ (.I(_04232_),
    .ZN(_00995_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08647_ (.I(\u_cpu.cpu.genblk3.csr.timer_irq_r ),
    .ZN(_04233_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08648_ (.A1(_02263_),
    .A2(_02598_),
    .Z(_04234_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _08649_ (.A1(\u_cpu.cpu.genblk3.csr.mie_mtie ),
    .A2(\u_cpu.cpu.genblk3.csr.mstatus_mie ),
    .A3(\u_cpu.cpu.genblk3.csr.i_mtip ),
    .A4(_04234_),
    .ZN(_04235_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08650_ (.A1(_04233_),
    .A2(_04234_),
    .B(_04235_),
    .ZN(_00996_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08651_ (.A1(_02754_),
    .A2(_02782_),
    .ZN(_04236_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08652_ (.I(_04236_),
    .Z(_04237_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08653_ (.A1(\u_cpu.rf_ram.memory[32][0] ),
    .A2(_04237_),
    .ZN(_04238_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08654_ (.A1(_03691_),
    .A2(_04237_),
    .B(_04238_),
    .ZN(_00997_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08655_ (.A1(\u_cpu.rf_ram.memory[32][1] ),
    .A2(_04237_),
    .ZN(_04239_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08656_ (.A1(_03695_),
    .A2(_04237_),
    .B(_04239_),
    .ZN(_00998_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08657_ (.A1(\u_cpu.rf_ram.memory[32][2] ),
    .A2(_04237_),
    .ZN(_04240_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08658_ (.A1(_03697_),
    .A2(_04237_),
    .B(_04240_),
    .ZN(_00999_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08659_ (.A1(\u_cpu.rf_ram.memory[32][3] ),
    .A2(_04237_),
    .ZN(_04241_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08660_ (.A1(_03699_),
    .A2(_04237_),
    .B(_04241_),
    .ZN(_01000_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08661_ (.A1(\u_cpu.rf_ram.memory[32][4] ),
    .A2(_04237_),
    .ZN(_04242_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08662_ (.A1(_03701_),
    .A2(_04237_),
    .B(_04242_),
    .ZN(_01001_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08663_ (.A1(\u_cpu.rf_ram.memory[32][5] ),
    .A2(_04237_),
    .ZN(_04243_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08664_ (.A1(_03703_),
    .A2(_04237_),
    .B(_04243_),
    .ZN(_01002_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08665_ (.A1(\u_cpu.rf_ram.memory[32][6] ),
    .A2(_04237_),
    .ZN(_04244_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08666_ (.A1(_03705_),
    .A2(_04237_),
    .B(_04244_),
    .ZN(_01003_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08667_ (.A1(\u_cpu.rf_ram.memory[32][7] ),
    .A2(_04237_),
    .ZN(_04245_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08668_ (.A1(_03707_),
    .A2(_04237_),
    .B(_04245_),
    .ZN(_01004_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08669_ (.A1(_02677_),
    .A2(_02870_),
    .ZN(_04246_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08670_ (.I(_04246_),
    .Z(_04247_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08671_ (.A1(\u_cpu.rf_ram.memory[31][0] ),
    .A2(_04247_),
    .ZN(_04248_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08672_ (.A1(_03691_),
    .A2(_04247_),
    .B(_04248_),
    .ZN(_01005_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08673_ (.A1(\u_cpu.rf_ram.memory[31][1] ),
    .A2(_04247_),
    .ZN(_04249_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08674_ (.A1(_03695_),
    .A2(_04247_),
    .B(_04249_),
    .ZN(_01006_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08675_ (.A1(\u_cpu.rf_ram.memory[31][2] ),
    .A2(_04247_),
    .ZN(_04250_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08676_ (.A1(_03697_),
    .A2(_04247_),
    .B(_04250_),
    .ZN(_01007_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08677_ (.A1(\u_cpu.rf_ram.memory[31][3] ),
    .A2(_04247_),
    .ZN(_04251_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08678_ (.A1(_03699_),
    .A2(_04247_),
    .B(_04251_),
    .ZN(_01008_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08679_ (.A1(\u_cpu.rf_ram.memory[31][4] ),
    .A2(_04247_),
    .ZN(_04252_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08680_ (.A1(_03701_),
    .A2(_04247_),
    .B(_04252_),
    .ZN(_01009_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08681_ (.A1(\u_cpu.rf_ram.memory[31][5] ),
    .A2(_04247_),
    .ZN(_04253_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08682_ (.A1(_03703_),
    .A2(_04247_),
    .B(_04253_),
    .ZN(_01010_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08683_ (.A1(\u_cpu.rf_ram.memory[31][6] ),
    .A2(_04247_),
    .ZN(_04254_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08684_ (.A1(_03705_),
    .A2(_04247_),
    .B(_04254_),
    .ZN(_01011_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08685_ (.A1(\u_cpu.rf_ram.memory[31][7] ),
    .A2(_04247_),
    .ZN(_04255_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08686_ (.A1(_03707_),
    .A2(_04247_),
    .B(_04255_),
    .ZN(_01012_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08687_ (.A1(\u_cpu.cpu.alu.cmp_r ),
    .A2(_02392_),
    .ZN(_04256_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08688_ (.A1(_02392_),
    .A2(_03646_),
    .B(_04256_),
    .ZN(_01013_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08689_ (.I(_02335_),
    .Z(_04257_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08690_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[2] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[3] ),
    .S(_04257_),
    .Z(_04258_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08691_ (.I(_04258_),
    .Z(_01014_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08692_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[3] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[4] ),
    .S(_04257_),
    .Z(_04259_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08693_ (.I(_04259_),
    .Z(_01015_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08694_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[4] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[5] ),
    .S(_04257_),
    .Z(_04260_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08695_ (.I(_04260_),
    .Z(_01016_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08696_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[5] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[6] ),
    .S(_04257_),
    .Z(_04261_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08697_ (.I(_04261_),
    .Z(_01017_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08698_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[6] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[7] ),
    .S(_04257_),
    .Z(_04262_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08699_ (.I(_04262_),
    .Z(_01018_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08700_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[7] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[8] ),
    .S(_04257_),
    .Z(_04263_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08701_ (.I(_04263_),
    .Z(_01019_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08702_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[8] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[9] ),
    .S(_04257_),
    .Z(_04264_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08703_ (.I(_04264_),
    .Z(_01020_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08704_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[9] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[10] ),
    .S(_04257_),
    .Z(_04265_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08705_ (.I(_04265_),
    .Z(_01021_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08706_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[10] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[11] ),
    .S(_04257_),
    .Z(_04266_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08707_ (.I(_04266_),
    .Z(_01022_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08708_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[11] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[12] ),
    .S(_04257_),
    .Z(_04267_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08709_ (.I(_04267_),
    .Z(_01023_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08710_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[12] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[13] ),
    .S(_04257_),
    .Z(_04268_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08711_ (.I(_04268_),
    .Z(_01024_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08712_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[13] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[14] ),
    .S(_04257_),
    .Z(_04269_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08713_ (.I(_04269_),
    .Z(_01025_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08714_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[14] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[15] ),
    .S(_04257_),
    .Z(_04270_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08715_ (.I(_04270_),
    .Z(_01026_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08716_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[15] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[16] ),
    .S(_04257_),
    .Z(_04271_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08717_ (.I(_04271_),
    .Z(_01027_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08718_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[16] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[17] ),
    .S(_04257_),
    .Z(_04272_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08719_ (.I(_04272_),
    .Z(_01028_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08720_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[17] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[18] ),
    .S(_04257_),
    .Z(_04273_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08721_ (.I(_04273_),
    .Z(_01029_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08722_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[18] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[19] ),
    .S(_02335_),
    .Z(_04274_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08723_ (.I(_04274_),
    .Z(_01030_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08724_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[19] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[20] ),
    .S(_02335_),
    .Z(_04275_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08725_ (.I(_04275_),
    .Z(_01031_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08726_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[20] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[21] ),
    .S(_02335_),
    .Z(_04276_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08727_ (.I(_04276_),
    .Z(_01032_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08728_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[21] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[22] ),
    .S(_02335_),
    .Z(_04277_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08729_ (.I(_04277_),
    .Z(_01033_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08730_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[22] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[23] ),
    .S(_02335_),
    .Z(_04278_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08731_ (.I(_04278_),
    .Z(_01034_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08732_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[23] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[24] ),
    .S(_02335_),
    .Z(_04279_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08733_ (.I(_04279_),
    .Z(_01035_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08734_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[24] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[25] ),
    .S(_02335_),
    .Z(_04280_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08735_ (.I(_04280_),
    .Z(_01036_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08736_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[25] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[26] ),
    .S(_02335_),
    .Z(_04281_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08737_ (.I(_04281_),
    .Z(_01037_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08738_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[26] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[27] ),
    .S(_02335_),
    .Z(_04282_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08739_ (.I(_04282_),
    .Z(_01038_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08740_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[27] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[28] ),
    .S(_02335_),
    .Z(_04283_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08741_ (.I(_04283_),
    .Z(_01039_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08742_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[28] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[29] ),
    .S(_02335_),
    .Z(_04284_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08743_ (.I(_04284_),
    .Z(_01040_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08744_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[29] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[30] ),
    .S(_02335_),
    .Z(_04285_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08745_ (.I(_04285_),
    .Z(_01041_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08746_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[30] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[31] ),
    .S(_02335_),
    .Z(_04286_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08747_ (.I(_04286_),
    .Z(_01042_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08748_ (.A1(_02590_),
    .A2(_02592_),
    .B(_02598_),
    .ZN(_04287_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08749_ (.A1(_02590_),
    .A2(_02592_),
    .B(_04287_),
    .ZN(_04288_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08750_ (.A1(\u_cpu.cpu.bufreg.i_sh_signed ),
    .A2(\u_arbiter.i_wb_cpu_dbus_adr[31] ),
    .A3(_02598_),
    .ZN(_04289_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08751_ (.A1(_04288_),
    .A2(_04289_),
    .ZN(_04290_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08752_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[31] ),
    .I1(_04290_),
    .S(_02335_),
    .Z(_04291_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08753_ (.I(_04291_),
    .Z(_01043_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08754_ (.A1(\u_cpu.cpu.state.o_cnt_r[1] ),
    .A2(\u_cpu.cpu.state.o_cnt_r[0] ),
    .B(_02292_),
    .C(_02914_),
    .ZN(_04292_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08755_ (.A1(_02596_),
    .A2(_02914_),
    .B(_04292_),
    .ZN(_04293_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08756_ (.A1(_02355_),
    .A2(_04293_),
    .ZN(_04294_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08757_ (.A1(_02412_),
    .A2(_04293_),
    .B(_04294_),
    .ZN(_01044_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08758_ (.A1(\u_arbiter.i_wb_cpu_dbus_adr[2] ),
    .A2(_02598_),
    .ZN(_04295_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08759_ (.A1(_04288_),
    .A2(_04295_),
    .ZN(_04296_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08760_ (.I0(_02355_),
    .I1(_04296_),
    .S(_04293_),
    .Z(_04297_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08761_ (.I(_04297_),
    .Z(_01045_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08762_ (.A1(_02677_),
    .A2(_02766_),
    .ZN(_04298_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08763_ (.I(_04298_),
    .Z(_04299_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08764_ (.A1(\u_cpu.rf_ram.memory[30][0] ),
    .A2(_04299_),
    .ZN(_04300_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08765_ (.A1(_03691_),
    .A2(_04299_),
    .B(_04300_),
    .ZN(_01046_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08766_ (.A1(\u_cpu.rf_ram.memory[30][1] ),
    .A2(_04299_),
    .ZN(_04301_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08767_ (.A1(_03695_),
    .A2(_04299_),
    .B(_04301_),
    .ZN(_01047_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08768_ (.A1(\u_cpu.rf_ram.memory[30][2] ),
    .A2(_04299_),
    .ZN(_04302_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08769_ (.A1(_03697_),
    .A2(_04299_),
    .B(_04302_),
    .ZN(_01048_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08770_ (.A1(\u_cpu.rf_ram.memory[30][3] ),
    .A2(_04299_),
    .ZN(_04303_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08771_ (.A1(_03699_),
    .A2(_04299_),
    .B(_04303_),
    .ZN(_01049_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08772_ (.A1(\u_cpu.rf_ram.memory[30][4] ),
    .A2(_04299_),
    .ZN(_04304_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08773_ (.A1(_03701_),
    .A2(_04299_),
    .B(_04304_),
    .ZN(_01050_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08774_ (.A1(\u_cpu.rf_ram.memory[30][5] ),
    .A2(_04299_),
    .ZN(_04305_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08775_ (.A1(_03703_),
    .A2(_04299_),
    .B(_04305_),
    .ZN(_01051_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08776_ (.A1(\u_cpu.rf_ram.memory[30][6] ),
    .A2(_04299_),
    .ZN(_04306_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08777_ (.A1(_03705_),
    .A2(_04299_),
    .B(_04306_),
    .ZN(_01052_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08778_ (.A1(\u_cpu.rf_ram.memory[30][7] ),
    .A2(_04299_),
    .ZN(_04307_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08779_ (.A1(_03707_),
    .A2(_04299_),
    .B(_04307_),
    .ZN(_01053_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08780_ (.A1(_02259_),
    .A2(_02598_),
    .B(_02395_),
    .ZN(_04308_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08781_ (.I(_04308_),
    .Z(_04309_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08782_ (.A1(_02395_),
    .A2(_02599_),
    .ZN(_04310_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08783_ (.I(_04310_),
    .Z(_04311_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08784_ (.A1(\u_arbiter.i_wb_cpu_ibus_adr[0] ),
    .A2(_04309_),
    .B1(_04311_),
    .B2(\u_arbiter.i_wb_cpu_ibus_adr[1] ),
    .ZN(_04312_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _08785_ (.I(_04312_),
    .ZN(_01054_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08786_ (.A1(\u_arbiter.i_wb_cpu_ibus_adr[1] ),
    .A2(_04309_),
    .B1(_04311_),
    .B2(\u_cpu.cpu.ctrl.o_ibus_adr[2] ),
    .ZN(_04313_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _08787_ (.I(_04313_),
    .ZN(_01055_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08788_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[2] ),
    .A2(_04309_),
    .B1(_04311_),
    .B2(\u_cpu.cpu.ctrl.o_ibus_adr[3] ),
    .ZN(_04314_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _08789_ (.I(_04314_),
    .ZN(_01056_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08790_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[3] ),
    .A2(_04309_),
    .B1(_04311_),
    .B2(\u_cpu.cpu.ctrl.o_ibus_adr[4] ),
    .ZN(_04315_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _08791_ (.I(_04315_),
    .ZN(_01057_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08792_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[4] ),
    .A2(_04309_),
    .B1(_04311_),
    .B2(\u_cpu.cpu.ctrl.o_ibus_adr[5] ),
    .ZN(_04316_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _08793_ (.I(_04316_),
    .ZN(_01058_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08794_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[5] ),
    .A2(_04309_),
    .B1(_04311_),
    .B2(\u_cpu.cpu.ctrl.o_ibus_adr[6] ),
    .ZN(_04317_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _08795_ (.I(_04317_),
    .ZN(_01059_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08796_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[6] ),
    .A2(_04309_),
    .B1(_04311_),
    .B2(\u_cpu.cpu.ctrl.o_ibus_adr[7] ),
    .ZN(_04318_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _08797_ (.I(_04318_),
    .ZN(_01060_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08798_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[7] ),
    .A2(_04309_),
    .B1(_04311_),
    .B2(\u_cpu.cpu.ctrl.o_ibus_adr[8] ),
    .ZN(_04319_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _08799_ (.I(_04319_),
    .ZN(_01061_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08800_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[8] ),
    .A2(_04309_),
    .B1(_04311_),
    .B2(\u_cpu.cpu.ctrl.o_ibus_adr[9] ),
    .ZN(_04320_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _08801_ (.I(_04320_),
    .ZN(_01062_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08802_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[9] ),
    .A2(_04309_),
    .B1(_04311_),
    .B2(\u_cpu.cpu.ctrl.o_ibus_adr[10] ),
    .ZN(_04321_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _08803_ (.I(_04321_),
    .ZN(_01063_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08804_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[10] ),
    .A2(_04309_),
    .B1(_04311_),
    .B2(\u_cpu.cpu.ctrl.o_ibus_adr[11] ),
    .ZN(_04322_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _08805_ (.I(_04322_),
    .ZN(_01064_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08806_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[11] ),
    .A2(_04309_),
    .B1(_04311_),
    .B2(\u_cpu.cpu.ctrl.o_ibus_adr[12] ),
    .ZN(_04323_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _08807_ (.I(_04323_),
    .ZN(_01065_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08808_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[12] ),
    .A2(_04309_),
    .B1(_04311_),
    .B2(\u_cpu.cpu.ctrl.o_ibus_adr[13] ),
    .ZN(_04324_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _08809_ (.I(_04324_),
    .ZN(_01066_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08810_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[13] ),
    .A2(_04309_),
    .B1(_04311_),
    .B2(\u_cpu.cpu.ctrl.o_ibus_adr[14] ),
    .ZN(_04325_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _08811_ (.I(_04325_),
    .ZN(_01067_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08812_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[14] ),
    .A2(_04309_),
    .B1(_04311_),
    .B2(\u_cpu.cpu.ctrl.o_ibus_adr[15] ),
    .ZN(_04326_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _08813_ (.I(_04326_),
    .ZN(_01068_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08814_ (.I(_04308_),
    .Z(_04327_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08815_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[15] ),
    .A2(_04327_),
    .B1(_04311_),
    .B2(\u_cpu.cpu.ctrl.o_ibus_adr[16] ),
    .ZN(_04328_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _08816_ (.I(_04328_),
    .ZN(_01069_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08817_ (.I(_04310_),
    .Z(_04329_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08818_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[16] ),
    .A2(_04327_),
    .B1(_04329_),
    .B2(\u_cpu.cpu.ctrl.o_ibus_adr[17] ),
    .ZN(_04330_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _08819_ (.I(_04330_),
    .ZN(_01070_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08820_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[17] ),
    .A2(_04327_),
    .B1(_04329_),
    .B2(\u_cpu.cpu.ctrl.o_ibus_adr[18] ),
    .ZN(_04331_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _08821_ (.I(_04331_),
    .ZN(_01071_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08822_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[18] ),
    .A2(_04327_),
    .B1(_04329_),
    .B2(\u_cpu.cpu.ctrl.o_ibus_adr[19] ),
    .ZN(_04332_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _08823_ (.I(_04332_),
    .ZN(_01072_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08824_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[19] ),
    .A2(_04327_),
    .B1(_04329_),
    .B2(\u_cpu.cpu.ctrl.o_ibus_adr[20] ),
    .ZN(_04333_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _08825_ (.I(_04333_),
    .ZN(_01073_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08826_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[20] ),
    .A2(_04327_),
    .B1(_04329_),
    .B2(\u_cpu.cpu.ctrl.o_ibus_adr[21] ),
    .ZN(_04334_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _08827_ (.I(_04334_),
    .ZN(_01074_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08828_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[21] ),
    .A2(_04327_),
    .B1(_04329_),
    .B2(\u_cpu.cpu.ctrl.o_ibus_adr[22] ),
    .ZN(_04335_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _08829_ (.I(_04335_),
    .ZN(_01075_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08830_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[22] ),
    .A2(_04327_),
    .B1(_04329_),
    .B2(\u_cpu.cpu.ctrl.o_ibus_adr[23] ),
    .ZN(_04336_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _08831_ (.I(_04336_),
    .ZN(_01076_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08832_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[23] ),
    .A2(_04327_),
    .B1(_04329_),
    .B2(\u_cpu.cpu.ctrl.o_ibus_adr[24] ),
    .ZN(_04337_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _08833_ (.I(_04337_),
    .ZN(_01077_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08834_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[24] ),
    .A2(_04327_),
    .B1(_04329_),
    .B2(\u_cpu.cpu.ctrl.o_ibus_adr[25] ),
    .ZN(_04338_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _08835_ (.I(_04338_),
    .ZN(_01078_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08836_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[25] ),
    .A2(_04327_),
    .B1(_04329_),
    .B2(\u_cpu.cpu.ctrl.o_ibus_adr[26] ),
    .ZN(_04339_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _08837_ (.I(_04339_),
    .ZN(_01079_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08838_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[26] ),
    .A2(_04327_),
    .B1(_04329_),
    .B2(\u_cpu.cpu.ctrl.o_ibus_adr[27] ),
    .ZN(_04340_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _08839_ (.I(_04340_),
    .ZN(_01080_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08840_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[27] ),
    .A2(_04327_),
    .B1(_04329_),
    .B2(\u_cpu.cpu.ctrl.o_ibus_adr[28] ),
    .ZN(_04341_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _08841_ (.I(_04341_),
    .ZN(_01081_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08842_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[28] ),
    .A2(_04327_),
    .B1(_04329_),
    .B2(\u_cpu.cpu.ctrl.o_ibus_adr[29] ),
    .ZN(_04342_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _08843_ (.I(_04342_),
    .ZN(_01082_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08844_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[29] ),
    .A2(_04327_),
    .B1(_04329_),
    .B2(\u_cpu.cpu.ctrl.o_ibus_adr[30] ),
    .ZN(_04343_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _08845_ (.I(_04343_),
    .ZN(_01083_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08846_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[30] ),
    .A2(_04327_),
    .B1(_04329_),
    .B2(\u_cpu.cpu.ctrl.o_ibus_adr[31] ),
    .ZN(_04344_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _08847_ (.I(_04344_),
    .ZN(_01084_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08848_ (.I0(_02363_),
    .I1(_02341_),
    .S(\u_cpu.cpu.ctrl.i_jump ),
    .Z(_04345_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08849_ (.A1(_02276_),
    .A2(_02334_),
    .B(_01451_),
    .ZN(_04346_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08850_ (.A1(_01451_),
    .A2(_04345_),
    .B(_04346_),
    .ZN(_04347_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08851_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[31] ),
    .A2(_04308_),
    .B1(_04329_),
    .B2(_04347_),
    .ZN(_04348_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _08852_ (.I(_04348_),
    .ZN(_01085_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _08853_ (.A1(\u_cpu.cpu.immdec.imm11_7[2] ),
    .A2(_02624_),
    .A3(_02729_),
    .ZN(_04349_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08854_ (.A1(_02803_),
    .A2(_04349_),
    .ZN(_04350_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08855_ (.I(_04350_),
    .Z(_04351_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08856_ (.A1(\u_cpu.rf_ram.memory[109][0] ),
    .A2(_04351_),
    .ZN(_04352_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08857_ (.A1(_03691_),
    .A2(_04351_),
    .B(_04352_),
    .ZN(_01086_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08858_ (.A1(\u_cpu.rf_ram.memory[109][1] ),
    .A2(_04351_),
    .ZN(_04353_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08859_ (.A1(_03695_),
    .A2(_04351_),
    .B(_04353_),
    .ZN(_01087_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08860_ (.A1(\u_cpu.rf_ram.memory[109][2] ),
    .A2(_04351_),
    .ZN(_04354_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08861_ (.A1(_03697_),
    .A2(_04351_),
    .B(_04354_),
    .ZN(_01088_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08862_ (.A1(\u_cpu.rf_ram.memory[109][3] ),
    .A2(_04351_),
    .ZN(_04355_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08863_ (.A1(_03699_),
    .A2(_04351_),
    .B(_04355_),
    .ZN(_01089_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08864_ (.A1(\u_cpu.rf_ram.memory[109][4] ),
    .A2(_04351_),
    .ZN(_04356_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08865_ (.A1(_03701_),
    .A2(_04351_),
    .B(_04356_),
    .ZN(_01090_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08866_ (.A1(\u_cpu.rf_ram.memory[109][5] ),
    .A2(_04351_),
    .ZN(_04357_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08867_ (.A1(_03703_),
    .A2(_04351_),
    .B(_04357_),
    .ZN(_01091_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08868_ (.A1(\u_cpu.rf_ram.memory[109][6] ),
    .A2(_04351_),
    .ZN(_04358_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08869_ (.A1(_03705_),
    .A2(_04351_),
    .B(_04358_),
    .ZN(_01092_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08870_ (.A1(\u_cpu.rf_ram.memory[109][7] ),
    .A2(_04351_),
    .ZN(_04359_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08871_ (.A1(_03707_),
    .A2(_04351_),
    .B(_04359_),
    .ZN(_01093_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08872_ (.A1(_02731_),
    .A2(_02825_),
    .Z(_04360_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08873_ (.I(_04360_),
    .Z(_04361_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08874_ (.A1(\u_cpu.rf_ram.memory[3][0] ),
    .A2(_04361_),
    .ZN(_04362_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08875_ (.A1(_02632_),
    .A2(_04361_),
    .B(_04362_),
    .ZN(_01094_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08876_ (.A1(\u_cpu.rf_ram.memory[3][1] ),
    .A2(_04361_),
    .ZN(_04363_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08877_ (.A1(_02637_),
    .A2(_04361_),
    .B(_04363_),
    .ZN(_01095_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08878_ (.A1(\u_cpu.rf_ram.memory[3][2] ),
    .A2(_04361_),
    .ZN(_04364_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08879_ (.A1(_02642_),
    .A2(_04361_),
    .B(_04364_),
    .ZN(_01096_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08880_ (.A1(\u_cpu.rf_ram.memory[3][3] ),
    .A2(_04361_),
    .ZN(_04365_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08881_ (.A1(_02647_),
    .A2(_04361_),
    .B(_04365_),
    .ZN(_01097_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08882_ (.A1(\u_cpu.rf_ram.memory[3][4] ),
    .A2(_04361_),
    .ZN(_04366_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08883_ (.A1(_02652_),
    .A2(_04361_),
    .B(_04366_),
    .ZN(_01098_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08884_ (.A1(\u_cpu.rf_ram.memory[3][5] ),
    .A2(_04361_),
    .ZN(_04367_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08885_ (.A1(_02657_),
    .A2(_04361_),
    .B(_04367_),
    .ZN(_01099_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08886_ (.A1(\u_cpu.rf_ram.memory[3][6] ),
    .A2(_04361_),
    .ZN(_04368_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08887_ (.A1(_02662_),
    .A2(_04361_),
    .B(_04368_),
    .ZN(_01100_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08888_ (.A1(\u_cpu.rf_ram.memory[3][7] ),
    .A2(_04361_),
    .ZN(_04369_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08889_ (.A1(_02667_),
    .A2(_04361_),
    .B(_04369_),
    .ZN(_01101_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08890_ (.A1(_02619_),
    .A2(_02731_),
    .Z(_04370_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08891_ (.I(_04370_),
    .Z(_04371_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08892_ (.A1(\u_cpu.rf_ram.memory[2][0] ),
    .A2(_04371_),
    .ZN(_04372_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08893_ (.A1(_02632_),
    .A2(_04371_),
    .B(_04372_),
    .ZN(_01102_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08894_ (.A1(\u_cpu.rf_ram.memory[2][1] ),
    .A2(_04371_),
    .ZN(_04373_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08895_ (.A1(_02637_),
    .A2(_04371_),
    .B(_04373_),
    .ZN(_01103_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08896_ (.A1(\u_cpu.rf_ram.memory[2][2] ),
    .A2(_04371_),
    .ZN(_04374_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08897_ (.A1(_02642_),
    .A2(_04371_),
    .B(_04374_),
    .ZN(_01104_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08898_ (.A1(\u_cpu.rf_ram.memory[2][3] ),
    .A2(_04371_),
    .ZN(_04375_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08899_ (.A1(_02647_),
    .A2(_04371_),
    .B(_04375_),
    .ZN(_01105_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08900_ (.A1(\u_cpu.rf_ram.memory[2][4] ),
    .A2(_04371_),
    .ZN(_04376_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08901_ (.A1(_02652_),
    .A2(_04371_),
    .B(_04376_),
    .ZN(_01106_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08902_ (.A1(\u_cpu.rf_ram.memory[2][5] ),
    .A2(_04371_),
    .ZN(_04377_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08903_ (.A1(_02657_),
    .A2(_04371_),
    .B(_04377_),
    .ZN(_01107_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08904_ (.A1(\u_cpu.rf_ram.memory[2][6] ),
    .A2(_04371_),
    .ZN(_04378_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08905_ (.A1(_02662_),
    .A2(_04371_),
    .B(_04378_),
    .ZN(_01108_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08906_ (.A1(\u_cpu.rf_ram.memory[2][7] ),
    .A2(_04371_),
    .ZN(_04379_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08907_ (.A1(_02667_),
    .A2(_04371_),
    .B(_04379_),
    .ZN(_01109_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08908_ (.A1(_02626_),
    .A2(_02803_),
    .ZN(_04380_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08909_ (.I(_04380_),
    .Z(_04381_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08910_ (.A1(\u_cpu.rf_ram.memory[93][0] ),
    .A2(_04381_),
    .ZN(_04382_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08911_ (.A1(_03691_),
    .A2(_04381_),
    .B(_04382_),
    .ZN(_01110_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08912_ (.A1(\u_cpu.rf_ram.memory[93][1] ),
    .A2(_04381_),
    .ZN(_04383_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08913_ (.A1(_03695_),
    .A2(_04381_),
    .B(_04383_),
    .ZN(_01111_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08914_ (.A1(\u_cpu.rf_ram.memory[93][2] ),
    .A2(_04381_),
    .ZN(_04384_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08915_ (.A1(_03697_),
    .A2(_04381_),
    .B(_04384_),
    .ZN(_01112_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08916_ (.A1(\u_cpu.rf_ram.memory[93][3] ),
    .A2(_04381_),
    .ZN(_04385_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08917_ (.A1(_03699_),
    .A2(_04381_),
    .B(_04385_),
    .ZN(_01113_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08918_ (.A1(\u_cpu.rf_ram.memory[93][4] ),
    .A2(_04381_),
    .ZN(_04386_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08919_ (.A1(_03701_),
    .A2(_04381_),
    .B(_04386_),
    .ZN(_01114_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08920_ (.A1(\u_cpu.rf_ram.memory[93][5] ),
    .A2(_04381_),
    .ZN(_04387_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08921_ (.A1(_03703_),
    .A2(_04381_),
    .B(_04387_),
    .ZN(_01115_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08922_ (.A1(\u_cpu.rf_ram.memory[93][6] ),
    .A2(_04381_),
    .ZN(_04388_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08923_ (.A1(_03705_),
    .A2(_04381_),
    .B(_04388_),
    .ZN(_01116_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08924_ (.A1(\u_cpu.rf_ram.memory[93][7] ),
    .A2(_04381_),
    .ZN(_04389_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08925_ (.A1(_03707_),
    .A2(_04381_),
    .B(_04389_),
    .ZN(_01117_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08926_ (.A1(_02392_),
    .A2(_02604_),
    .ZN(_04390_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08927_ (.A1(_03955_),
    .A2(_04390_),
    .ZN(_04391_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08928_ (.A1(\u_cpu.cpu.immdec.imm11_7[1] ),
    .A2(_03897_),
    .B(_04391_),
    .ZN(_04392_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08929_ (.A1(_02264_),
    .A2(_04391_),
    .B1(_04392_),
    .B2(_04160_),
    .ZN(_01118_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _08930_ (.A1(_03932_),
    .A2(_03939_),
    .A3(_03948_),
    .A4(_03962_),
    .ZN(_04393_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _08931_ (.A1(_03932_),
    .A2(_03975_),
    .B1(_03988_),
    .B2(_03944_),
    .C(_04188_),
    .ZN(_04394_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _08932_ (.A1(_03928_),
    .A2(_04188_),
    .B1(_04190_),
    .B2(_04394_),
    .C(_03969_),
    .ZN(_04395_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08933_ (.A1(_03910_),
    .A2(_04395_),
    .B(_03965_),
    .ZN(_04396_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08934_ (.A1(_03944_),
    .A2(_03908_),
    .B1(_03909_),
    .B2(_03932_),
    .ZN(_04397_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08935_ (.A1(_04393_),
    .A2(_04396_),
    .B1(_04397_),
    .B2(_03910_),
    .ZN(_04398_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08936_ (.A1(_03956_),
    .A2(_04398_),
    .ZN(_04399_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08937_ (.A1(\u_cpu.cpu.immdec.imm11_7[1] ),
    .A2(_04390_),
    .ZN(_04400_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08938_ (.A1(_02728_),
    .A2(_04390_),
    .B(_04400_),
    .ZN(_04401_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08939_ (.A1(_03932_),
    .A2(_04009_),
    .B1(_04401_),
    .B2(_03897_),
    .ZN(_04402_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08940_ (.A1(_04399_),
    .A2(_04402_),
    .ZN(_01119_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08941_ (.A1(_03986_),
    .A2(_03949_),
    .B(_03965_),
    .ZN(_04403_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08942_ (.A1(_03924_),
    .A2(_04403_),
    .ZN(_04404_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08943_ (.A1(_03924_),
    .A2(_03977_),
    .A3(_03985_),
    .ZN(_04405_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08944_ (.A1(_03945_),
    .A2(_03988_),
    .B(_04188_),
    .ZN(_04406_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08945_ (.A1(_04405_),
    .A2(_04406_),
    .B(_04179_),
    .ZN(_04407_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08946_ (.A1(_03940_),
    .A2(_03910_),
    .ZN(_04408_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _08947_ (.A1(_03958_),
    .A2(_03947_),
    .A3(_04031_),
    .B1(_03962_),
    .B2(_04408_),
    .ZN(_04409_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _08948_ (.A1(_03896_),
    .A2(_04407_),
    .A3(_04409_),
    .ZN(_04410_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08949_ (.A1(_02728_),
    .A2(_04390_),
    .ZN(_04411_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08950_ (.A1(\u_cpu.cpu.immdec.imm11_7[3] ),
    .A2(_04390_),
    .B(_04411_),
    .C(_03955_),
    .ZN(_04412_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08951_ (.A1(_04404_),
    .A2(_04410_),
    .B(_04412_),
    .ZN(_01120_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _08952_ (.A1(\u_cpu.cpu.immdec.imm11_7[4] ),
    .A2(_02392_),
    .A3(_02604_),
    .ZN(_04413_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08953_ (.A1(\u_cpu.cpu.immdec.imm11_7[3] ),
    .A2(_04390_),
    .B(_03897_),
    .ZN(_04414_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08954_ (.A1(_03903_),
    .A2(_03918_),
    .B(_04031_),
    .ZN(_04415_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08955_ (.A1(_04403_),
    .A2(_04415_),
    .B(_03923_),
    .ZN(_04416_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _08956_ (.A1(_03947_),
    .A2(_04031_),
    .B1(_03969_),
    .B2(_03970_),
    .C(_04416_),
    .ZN(_04417_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08957_ (.A1(_03956_),
    .A2(_04417_),
    .ZN(_04418_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08958_ (.A1(_04413_),
    .A2(_04414_),
    .B(_04418_),
    .ZN(_01121_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08959_ (.A1(_03901_),
    .A2(_03919_),
    .ZN(_04419_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08960_ (.A1(_04024_),
    .A2(_04419_),
    .B(_03948_),
    .C(_04031_),
    .ZN(_04420_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08961_ (.A1(_03965_),
    .A2(_03962_),
    .A3(_04420_),
    .ZN(_04421_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08962_ (.A1(_03956_),
    .A2(_03922_),
    .A3(_04421_),
    .ZN(_04422_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08963_ (.A1(\u_cpu.cpu.immdec.imm30_25[0] ),
    .A2(_03897_),
    .B(_04391_),
    .ZN(_04423_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08964_ (.A1(_02621_),
    .A2(_04391_),
    .B1(_04422_),
    .B2(_04423_),
    .ZN(_01122_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08965_ (.A1(_02695_),
    .A2(_04349_),
    .ZN(_04424_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08966_ (.I(_04424_),
    .Z(_04425_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08967_ (.A1(\u_cpu.rf_ram.memory[97][0] ),
    .A2(_04425_),
    .ZN(_04426_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08968_ (.A1(_03691_),
    .A2(_04425_),
    .B(_04426_),
    .ZN(_01123_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08969_ (.A1(\u_cpu.rf_ram.memory[97][1] ),
    .A2(_04425_),
    .ZN(_04427_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08970_ (.A1(_03695_),
    .A2(_04425_),
    .B(_04427_),
    .ZN(_01124_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08971_ (.A1(\u_cpu.rf_ram.memory[97][2] ),
    .A2(_04425_),
    .ZN(_04428_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08972_ (.A1(_03697_),
    .A2(_04425_),
    .B(_04428_),
    .ZN(_01125_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08973_ (.A1(\u_cpu.rf_ram.memory[97][3] ),
    .A2(_04425_),
    .ZN(_04429_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08974_ (.A1(_03699_),
    .A2(_04425_),
    .B(_04429_),
    .ZN(_01126_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08975_ (.A1(\u_cpu.rf_ram.memory[97][4] ),
    .A2(_04425_),
    .ZN(_04430_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08976_ (.A1(_03701_),
    .A2(_04425_),
    .B(_04430_),
    .ZN(_01127_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08977_ (.A1(\u_cpu.rf_ram.memory[97][5] ),
    .A2(_04425_),
    .ZN(_04431_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08978_ (.A1(_03703_),
    .A2(_04425_),
    .B(_04431_),
    .ZN(_01128_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08979_ (.A1(\u_cpu.rf_ram.memory[97][6] ),
    .A2(_04425_),
    .ZN(_04432_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08980_ (.A1(_03705_),
    .A2(_04425_),
    .B(_04432_),
    .ZN(_01129_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08981_ (.A1(\u_cpu.rf_ram.memory[97][7] ),
    .A2(_04425_),
    .ZN(_04433_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08982_ (.A1(_03707_),
    .A2(_04425_),
    .B(_04433_),
    .ZN(_01130_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08983_ (.I(_02631_),
    .Z(_04434_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08984_ (.A1(_02626_),
    .A2(_02766_),
    .ZN(_04435_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08985_ (.I(_04435_),
    .Z(_04436_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08986_ (.A1(\u_cpu.rf_ram.memory[94][0] ),
    .A2(_04436_),
    .ZN(_04437_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08987_ (.A1(_04434_),
    .A2(_04436_),
    .B(_04437_),
    .ZN(_01131_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08988_ (.I(_02636_),
    .Z(_04438_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08989_ (.A1(\u_cpu.rf_ram.memory[94][1] ),
    .A2(_04436_),
    .ZN(_04439_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08990_ (.A1(_04438_),
    .A2(_04436_),
    .B(_04439_),
    .ZN(_01132_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08991_ (.I(_02641_),
    .Z(_04440_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08992_ (.A1(\u_cpu.rf_ram.memory[94][2] ),
    .A2(_04436_),
    .ZN(_04441_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08993_ (.A1(_04440_),
    .A2(_04436_),
    .B(_04441_),
    .ZN(_01133_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08994_ (.I(_02646_),
    .Z(_04442_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08995_ (.A1(\u_cpu.rf_ram.memory[94][3] ),
    .A2(_04436_),
    .ZN(_04443_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08996_ (.A1(_04442_),
    .A2(_04436_),
    .B(_04443_),
    .ZN(_01134_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08997_ (.I(_02651_),
    .Z(_04444_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08998_ (.A1(\u_cpu.rf_ram.memory[94][4] ),
    .A2(_04436_),
    .ZN(_04445_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08999_ (.A1(_04444_),
    .A2(_04436_),
    .B(_04445_),
    .ZN(_01135_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09000_ (.I(_02656_),
    .Z(_04446_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09001_ (.A1(\u_cpu.rf_ram.memory[94][5] ),
    .A2(_04436_),
    .ZN(_04447_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09002_ (.A1(_04446_),
    .A2(_04436_),
    .B(_04447_),
    .ZN(_01136_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09003_ (.I(_02661_),
    .Z(_04448_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09004_ (.A1(\u_cpu.rf_ram.memory[94][6] ),
    .A2(_04436_),
    .ZN(_04449_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09005_ (.A1(_04448_),
    .A2(_04436_),
    .B(_04449_),
    .ZN(_01137_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09006_ (.I(_02666_),
    .Z(_04450_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09007_ (.A1(\u_cpu.rf_ram.memory[94][7] ),
    .A2(_04436_),
    .ZN(_04451_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09008_ (.A1(_04450_),
    .A2(_04436_),
    .B(_04451_),
    .ZN(_01138_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09009_ (.A1(_02626_),
    .A2(_02870_),
    .ZN(_04452_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09010_ (.I(_04452_),
    .Z(_04453_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09011_ (.A1(\u_cpu.rf_ram.memory[95][0] ),
    .A2(_04453_),
    .ZN(_04454_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09012_ (.A1(_04434_),
    .A2(_04453_),
    .B(_04454_),
    .ZN(_01139_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09013_ (.A1(\u_cpu.rf_ram.memory[95][1] ),
    .A2(_04453_),
    .ZN(_04455_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09014_ (.A1(_04438_),
    .A2(_04453_),
    .B(_04455_),
    .ZN(_01140_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09015_ (.A1(\u_cpu.rf_ram.memory[95][2] ),
    .A2(_04453_),
    .ZN(_04456_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09016_ (.A1(_04440_),
    .A2(_04453_),
    .B(_04456_),
    .ZN(_01141_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09017_ (.A1(\u_cpu.rf_ram.memory[95][3] ),
    .A2(_04453_),
    .ZN(_04457_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09018_ (.A1(_04442_),
    .A2(_04453_),
    .B(_04457_),
    .ZN(_01142_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09019_ (.A1(\u_cpu.rf_ram.memory[95][4] ),
    .A2(_04453_),
    .ZN(_04458_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09020_ (.A1(_04444_),
    .A2(_04453_),
    .B(_04458_),
    .ZN(_01143_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09021_ (.A1(\u_cpu.rf_ram.memory[95][5] ),
    .A2(_04453_),
    .ZN(_04459_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09022_ (.A1(_04446_),
    .A2(_04453_),
    .B(_04459_),
    .ZN(_01144_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09023_ (.A1(\u_cpu.rf_ram.memory[95][6] ),
    .A2(_04453_),
    .ZN(_04460_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09024_ (.A1(_04448_),
    .A2(_04453_),
    .B(_04460_),
    .ZN(_01145_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09025_ (.A1(\u_cpu.rf_ram.memory[95][7] ),
    .A2(_04453_),
    .ZN(_04461_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09026_ (.A1(_04450_),
    .A2(_04453_),
    .B(_04461_),
    .ZN(_01146_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09027_ (.A1(_02754_),
    .A2(_04349_),
    .ZN(_04462_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09028_ (.I(_04462_),
    .Z(_04463_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09029_ (.A1(\u_cpu.rf_ram.memory[96][0] ),
    .A2(_04463_),
    .ZN(_04464_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09030_ (.A1(_04434_),
    .A2(_04463_),
    .B(_04464_),
    .ZN(_01147_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09031_ (.A1(\u_cpu.rf_ram.memory[96][1] ),
    .A2(_04463_),
    .ZN(_04465_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09032_ (.A1(_04438_),
    .A2(_04463_),
    .B(_04465_),
    .ZN(_01148_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09033_ (.A1(\u_cpu.rf_ram.memory[96][2] ),
    .A2(_04463_),
    .ZN(_04466_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09034_ (.A1(_04440_),
    .A2(_04463_),
    .B(_04466_),
    .ZN(_01149_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09035_ (.A1(\u_cpu.rf_ram.memory[96][3] ),
    .A2(_04463_),
    .ZN(_04467_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09036_ (.A1(_04442_),
    .A2(_04463_),
    .B(_04467_),
    .ZN(_01150_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09037_ (.A1(\u_cpu.rf_ram.memory[96][4] ),
    .A2(_04463_),
    .ZN(_04468_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09038_ (.A1(_04444_),
    .A2(_04463_),
    .B(_04468_),
    .ZN(_01151_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09039_ (.A1(\u_cpu.rf_ram.memory[96][5] ),
    .A2(_04463_),
    .ZN(_04469_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09040_ (.A1(_04446_),
    .A2(_04463_),
    .B(_04469_),
    .ZN(_01152_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09041_ (.A1(\u_cpu.rf_ram.memory[96][6] ),
    .A2(_04463_),
    .ZN(_04470_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09042_ (.A1(_04448_),
    .A2(_04463_),
    .B(_04470_),
    .ZN(_01153_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09043_ (.A1(\u_cpu.rf_ram.memory[96][7] ),
    .A2(_04463_),
    .ZN(_04471_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09044_ (.A1(_04450_),
    .A2(_04463_),
    .B(_04471_),
    .ZN(_01154_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09045_ (.A1(\u_cpu.cpu.bufreg.i_sh_signed ),
    .A2(_03897_),
    .ZN(_04472_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09046_ (.A1(_04141_),
    .A2(_04472_),
    .ZN(_01155_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09047_ (.A1(\u_arbiter.i_wb_cpu_ibus_adr[1] ),
    .A2(\u_arbiter.i_wb_cpu_ack ),
    .A3(_02461_),
    .ZN(_04473_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09048_ (.A1(_02467_),
    .A2(_04473_),
    .Z(_04474_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09049_ (.A1(_02395_),
    .A2(_04474_),
    .ZN(_01156_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09050_ (.A1(_02677_),
    .A2(_02814_),
    .ZN(_04475_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09051_ (.I(_04475_),
    .Z(_04476_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09052_ (.A1(\u_cpu.rf_ram.memory[28][0] ),
    .A2(_04476_),
    .ZN(_04477_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09053_ (.A1(_04434_),
    .A2(_04476_),
    .B(_04477_),
    .ZN(_01157_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09054_ (.A1(\u_cpu.rf_ram.memory[28][1] ),
    .A2(_04476_),
    .ZN(_04478_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09055_ (.A1(_04438_),
    .A2(_04476_),
    .B(_04478_),
    .ZN(_01158_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09056_ (.A1(\u_cpu.rf_ram.memory[28][2] ),
    .A2(_04476_),
    .ZN(_04479_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09057_ (.A1(_04440_),
    .A2(_04476_),
    .B(_04479_),
    .ZN(_01159_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09058_ (.A1(\u_cpu.rf_ram.memory[28][3] ),
    .A2(_04476_),
    .ZN(_04480_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09059_ (.A1(_04442_),
    .A2(_04476_),
    .B(_04480_),
    .ZN(_01160_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09060_ (.A1(\u_cpu.rf_ram.memory[28][4] ),
    .A2(_04476_),
    .ZN(_04481_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09061_ (.A1(_04444_),
    .A2(_04476_),
    .B(_04481_),
    .ZN(_01161_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09062_ (.A1(\u_cpu.rf_ram.memory[28][5] ),
    .A2(_04476_),
    .ZN(_04482_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09063_ (.A1(_04446_),
    .A2(_04476_),
    .B(_04482_),
    .ZN(_01162_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09064_ (.A1(\u_cpu.rf_ram.memory[28][6] ),
    .A2(_04476_),
    .ZN(_04483_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09065_ (.A1(_04448_),
    .A2(_04476_),
    .B(_04483_),
    .ZN(_01163_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09066_ (.A1(\u_cpu.rf_ram.memory[28][7] ),
    .A2(_04476_),
    .ZN(_04484_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09067_ (.A1(_04450_),
    .A2(_04476_),
    .B(_04484_),
    .ZN(_01164_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09068_ (.I(_02910_),
    .Z(_04485_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09069_ (.I0(\u_arbiter.i_wb_cpu_rdt[16] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[0] ),
    .S(_04485_),
    .Z(_04486_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09070_ (.I(_04486_),
    .Z(_01165_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09071_ (.I0(\u_arbiter.i_wb_cpu_rdt[17] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[1] ),
    .S(_04485_),
    .Z(_04487_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09072_ (.I(_04487_),
    .Z(_01166_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09073_ (.I0(\u_arbiter.i_wb_cpu_rdt[18] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[2] ),
    .S(_04485_),
    .Z(_04488_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09074_ (.I(_04488_),
    .Z(_01167_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09075_ (.I0(\u_arbiter.i_wb_cpu_rdt[19] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[3] ),
    .S(_04485_),
    .Z(_04489_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09076_ (.I(_04489_),
    .Z(_01168_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09077_ (.I0(\u_arbiter.i_wb_cpu_rdt[20] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[4] ),
    .S(_04485_),
    .Z(_04490_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09078_ (.I(_04490_),
    .Z(_01169_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09079_ (.I0(\u_arbiter.i_wb_cpu_rdt[21] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[5] ),
    .S(_04485_),
    .Z(_04491_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09080_ (.I(_04491_),
    .Z(_01170_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09081_ (.I0(\u_arbiter.i_wb_cpu_rdt[22] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[6] ),
    .S(_04485_),
    .Z(_04492_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09082_ (.I(_04492_),
    .Z(_01171_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09083_ (.I0(\u_arbiter.i_wb_cpu_rdt[23] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[7] ),
    .S(_04485_),
    .Z(_04493_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09084_ (.I(_04493_),
    .Z(_01172_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09085_ (.I0(\u_arbiter.i_wb_cpu_rdt[24] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[8] ),
    .S(_04485_),
    .Z(_04494_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09086_ (.I(_04494_),
    .Z(_01173_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09087_ (.I0(\u_arbiter.i_wb_cpu_rdt[25] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[9] ),
    .S(_04485_),
    .Z(_04495_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09088_ (.I(_04495_),
    .Z(_01174_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09089_ (.I0(\u_arbiter.i_wb_cpu_rdt[26] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[10] ),
    .S(_04485_),
    .Z(_04496_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09090_ (.I(_04496_),
    .Z(_01175_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09091_ (.A1(\u_arbiter.i_wb_cpu_rdt[27] ),
    .A2(_04485_),
    .ZN(_04497_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09092_ (.A1(_03920_),
    .A2(_04485_),
    .B(_04497_),
    .ZN(_01176_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09093_ (.I0(\u_arbiter.i_wb_cpu_rdt[28] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[12] ),
    .S(_04485_),
    .Z(_04498_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09094_ (.I(_04498_),
    .Z(_01177_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09095_ (.I0(\u_arbiter.i_wb_cpu_rdt[29] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[13] ),
    .S(_04485_),
    .Z(_04499_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09096_ (.I(_04499_),
    .Z(_01178_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09097_ (.I0(\u_arbiter.i_wb_cpu_rdt[30] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[14] ),
    .S(_04485_),
    .Z(_04500_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09098_ (.I(_04500_),
    .Z(_01179_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09099_ (.I0(\u_arbiter.i_wb_cpu_rdt[31] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[15] ),
    .S(_02910_),
    .Z(_04501_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09100_ (.I(_04501_),
    .Z(_01180_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09101_ (.A1(_02675_),
    .A2(_04349_),
    .ZN(_04502_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09102_ (.I(_04502_),
    .Z(_04503_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09103_ (.A1(\u_cpu.rf_ram.memory[101][0] ),
    .A2(_04503_),
    .ZN(_04504_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09104_ (.A1(_04434_),
    .A2(_04503_),
    .B(_04504_),
    .ZN(_01181_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09105_ (.A1(\u_cpu.rf_ram.memory[101][1] ),
    .A2(_04503_),
    .ZN(_04505_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09106_ (.A1(_04438_),
    .A2(_04503_),
    .B(_04505_),
    .ZN(_01182_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09107_ (.A1(\u_cpu.rf_ram.memory[101][2] ),
    .A2(_04503_),
    .ZN(_04506_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09108_ (.A1(_04440_),
    .A2(_04503_),
    .B(_04506_),
    .ZN(_01183_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09109_ (.A1(\u_cpu.rf_ram.memory[101][3] ),
    .A2(_04503_),
    .ZN(_04507_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09110_ (.A1(_04442_),
    .A2(_04503_),
    .B(_04507_),
    .ZN(_01184_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09111_ (.A1(\u_cpu.rf_ram.memory[101][4] ),
    .A2(_04503_),
    .ZN(_04508_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09112_ (.A1(_04444_),
    .A2(_04503_),
    .B(_04508_),
    .ZN(_01185_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09113_ (.A1(\u_cpu.rf_ram.memory[101][5] ),
    .A2(_04503_),
    .ZN(_04509_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09114_ (.A1(_04446_),
    .A2(_04503_),
    .B(_04509_),
    .ZN(_01186_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09115_ (.A1(\u_cpu.rf_ram.memory[101][6] ),
    .A2(_04503_),
    .ZN(_04510_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09116_ (.A1(_04448_),
    .A2(_04503_),
    .B(_04510_),
    .ZN(_01187_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09117_ (.A1(\u_cpu.rf_ram.memory[101][7] ),
    .A2(_04503_),
    .ZN(_04511_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09118_ (.A1(_04450_),
    .A2(_04503_),
    .B(_04511_),
    .ZN(_01188_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09119_ (.A1(_03037_),
    .A2(_04349_),
    .ZN(_04512_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09120_ (.I(_04512_),
    .Z(_04513_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09121_ (.A1(\u_cpu.rf_ram.memory[102][0] ),
    .A2(_04513_),
    .ZN(_04514_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09122_ (.A1(_04434_),
    .A2(_04513_),
    .B(_04514_),
    .ZN(_01189_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09123_ (.A1(\u_cpu.rf_ram.memory[102][1] ),
    .A2(_04513_),
    .ZN(_04515_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09124_ (.A1(_04438_),
    .A2(_04513_),
    .B(_04515_),
    .ZN(_01190_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09125_ (.A1(\u_cpu.rf_ram.memory[102][2] ),
    .A2(_04513_),
    .ZN(_04516_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09126_ (.A1(_04440_),
    .A2(_04513_),
    .B(_04516_),
    .ZN(_01191_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09127_ (.A1(\u_cpu.rf_ram.memory[102][3] ),
    .A2(_04513_),
    .ZN(_04517_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09128_ (.A1(_04442_),
    .A2(_04513_),
    .B(_04517_),
    .ZN(_01192_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09129_ (.A1(\u_cpu.rf_ram.memory[102][4] ),
    .A2(_04513_),
    .ZN(_04518_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09130_ (.A1(_04444_),
    .A2(_04513_),
    .B(_04518_),
    .ZN(_01193_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09131_ (.A1(\u_cpu.rf_ram.memory[102][5] ),
    .A2(_04513_),
    .ZN(_04519_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09132_ (.A1(_04446_),
    .A2(_04513_),
    .B(_04519_),
    .ZN(_01194_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09133_ (.A1(\u_cpu.rf_ram.memory[102][6] ),
    .A2(_04513_),
    .ZN(_04520_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09134_ (.A1(_04448_),
    .A2(_04513_),
    .B(_04520_),
    .ZN(_01195_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09135_ (.A1(\u_cpu.rf_ram.memory[102][7] ),
    .A2(_04513_),
    .ZN(_04521_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09136_ (.A1(_04450_),
    .A2(_04513_),
    .B(_04521_),
    .ZN(_01196_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09137_ (.A1(_02743_),
    .A2(_04349_),
    .ZN(_04522_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09138_ (.I(_04522_),
    .Z(_04523_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09139_ (.A1(\u_cpu.rf_ram.memory[103][0] ),
    .A2(_04523_),
    .ZN(_04524_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09140_ (.A1(_04434_),
    .A2(_04523_),
    .B(_04524_),
    .ZN(_01197_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09141_ (.A1(\u_cpu.rf_ram.memory[103][1] ),
    .A2(_04523_),
    .ZN(_04525_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09142_ (.A1(_04438_),
    .A2(_04523_),
    .B(_04525_),
    .ZN(_01198_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09143_ (.A1(\u_cpu.rf_ram.memory[103][2] ),
    .A2(_04523_),
    .ZN(_04526_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09144_ (.A1(_04440_),
    .A2(_04523_),
    .B(_04526_),
    .ZN(_01199_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09145_ (.A1(\u_cpu.rf_ram.memory[103][3] ),
    .A2(_04523_),
    .ZN(_04527_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09146_ (.A1(_04442_),
    .A2(_04523_),
    .B(_04527_),
    .ZN(_01200_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09147_ (.A1(\u_cpu.rf_ram.memory[103][4] ),
    .A2(_04523_),
    .ZN(_04528_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09148_ (.A1(_04444_),
    .A2(_04523_),
    .B(_04528_),
    .ZN(_01201_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09149_ (.A1(\u_cpu.rf_ram.memory[103][5] ),
    .A2(_04523_),
    .ZN(_04529_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09150_ (.A1(_04446_),
    .A2(_04523_),
    .B(_04529_),
    .ZN(_01202_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09151_ (.A1(\u_cpu.rf_ram.memory[103][6] ),
    .A2(_04523_),
    .ZN(_04530_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09152_ (.A1(_04448_),
    .A2(_04523_),
    .B(_04530_),
    .ZN(_01203_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09153_ (.A1(\u_cpu.rf_ram.memory[103][7] ),
    .A2(_04523_),
    .ZN(_04531_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09154_ (.A1(_04450_),
    .A2(_04523_),
    .B(_04531_),
    .ZN(_01204_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09155_ (.A1(_02954_),
    .A2(_04349_),
    .ZN(_04532_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09156_ (.I(_04532_),
    .Z(_04533_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09157_ (.A1(\u_cpu.rf_ram.memory[104][0] ),
    .A2(_04533_),
    .ZN(_04534_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09158_ (.A1(_04434_),
    .A2(_04533_),
    .B(_04534_),
    .ZN(_01205_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09159_ (.A1(\u_cpu.rf_ram.memory[104][1] ),
    .A2(_04533_),
    .ZN(_04535_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09160_ (.A1(_04438_),
    .A2(_04533_),
    .B(_04535_),
    .ZN(_01206_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09161_ (.A1(\u_cpu.rf_ram.memory[104][2] ),
    .A2(_04533_),
    .ZN(_04536_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09162_ (.A1(_04440_),
    .A2(_04533_),
    .B(_04536_),
    .ZN(_01207_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09163_ (.A1(\u_cpu.rf_ram.memory[104][3] ),
    .A2(_04533_),
    .ZN(_04537_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09164_ (.A1(_04442_),
    .A2(_04533_),
    .B(_04537_),
    .ZN(_01208_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09165_ (.A1(\u_cpu.rf_ram.memory[104][4] ),
    .A2(_04533_),
    .ZN(_04538_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09166_ (.A1(_04444_),
    .A2(_04533_),
    .B(_04538_),
    .ZN(_01209_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09167_ (.A1(\u_cpu.rf_ram.memory[104][5] ),
    .A2(_04533_),
    .ZN(_04539_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09168_ (.A1(_04446_),
    .A2(_04533_),
    .B(_04539_),
    .ZN(_01210_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09169_ (.A1(\u_cpu.rf_ram.memory[104][6] ),
    .A2(_04533_),
    .ZN(_04540_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09170_ (.A1(_04448_),
    .A2(_04533_),
    .B(_04540_),
    .ZN(_01211_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09171_ (.A1(\u_cpu.rf_ram.memory[104][7] ),
    .A2(_04533_),
    .ZN(_04541_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09172_ (.A1(_04450_),
    .A2(_04533_),
    .B(_04541_),
    .ZN(_01212_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09173_ (.A1(_02825_),
    .A2(_04349_),
    .ZN(_04542_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09174_ (.I(_04542_),
    .Z(_04543_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09175_ (.A1(\u_cpu.rf_ram.memory[99][0] ),
    .A2(_04543_),
    .ZN(_04544_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09176_ (.A1(_04434_),
    .A2(_04543_),
    .B(_04544_),
    .ZN(_01213_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09177_ (.A1(\u_cpu.rf_ram.memory[99][1] ),
    .A2(_04543_),
    .ZN(_04545_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09178_ (.A1(_04438_),
    .A2(_04543_),
    .B(_04545_),
    .ZN(_01214_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09179_ (.A1(\u_cpu.rf_ram.memory[99][2] ),
    .A2(_04543_),
    .ZN(_04546_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09180_ (.A1(_04440_),
    .A2(_04543_),
    .B(_04546_),
    .ZN(_01215_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09181_ (.A1(\u_cpu.rf_ram.memory[99][3] ),
    .A2(_04543_),
    .ZN(_04547_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09182_ (.A1(_04442_),
    .A2(_04543_),
    .B(_04547_),
    .ZN(_01216_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09183_ (.A1(\u_cpu.rf_ram.memory[99][4] ),
    .A2(_04543_),
    .ZN(_04548_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09184_ (.A1(_04444_),
    .A2(_04543_),
    .B(_04548_),
    .ZN(_01217_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09185_ (.A1(\u_cpu.rf_ram.memory[99][5] ),
    .A2(_04543_),
    .ZN(_04549_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09186_ (.A1(_04446_),
    .A2(_04543_),
    .B(_04549_),
    .ZN(_01218_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09187_ (.A1(\u_cpu.rf_ram.memory[99][6] ),
    .A2(_04543_),
    .ZN(_04550_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09188_ (.A1(_04448_),
    .A2(_04543_),
    .B(_04550_),
    .ZN(_01219_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09189_ (.A1(\u_cpu.rf_ram.memory[99][7] ),
    .A2(_04543_),
    .ZN(_04551_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09190_ (.A1(_04450_),
    .A2(_04543_),
    .B(_04551_),
    .ZN(_01220_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09191_ (.A1(_02768_),
    .A2(_02870_),
    .ZN(_04552_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09192_ (.I(_04552_),
    .Z(_04553_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09193_ (.A1(\u_cpu.rf_ram.memory[79][0] ),
    .A2(_04553_),
    .ZN(_04554_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09194_ (.A1(_04434_),
    .A2(_04553_),
    .B(_04554_),
    .ZN(_01221_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09195_ (.A1(\u_cpu.rf_ram.memory[79][1] ),
    .A2(_04553_),
    .ZN(_04555_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09196_ (.A1(_04438_),
    .A2(_04553_),
    .B(_04555_),
    .ZN(_01222_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09197_ (.A1(\u_cpu.rf_ram.memory[79][2] ),
    .A2(_04553_),
    .ZN(_04556_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09198_ (.A1(_04440_),
    .A2(_04553_),
    .B(_04556_),
    .ZN(_01223_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09199_ (.A1(\u_cpu.rf_ram.memory[79][3] ),
    .A2(_04553_),
    .ZN(_04557_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09200_ (.A1(_04442_),
    .A2(_04553_),
    .B(_04557_),
    .ZN(_01224_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09201_ (.A1(\u_cpu.rf_ram.memory[79][4] ),
    .A2(_04553_),
    .ZN(_04558_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09202_ (.A1(_04444_),
    .A2(_04553_),
    .B(_04558_),
    .ZN(_01225_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09203_ (.A1(\u_cpu.rf_ram.memory[79][5] ),
    .A2(_04553_),
    .ZN(_04559_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09204_ (.A1(_04446_),
    .A2(_04553_),
    .B(_04559_),
    .ZN(_01226_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09205_ (.A1(\u_cpu.rf_ram.memory[79][6] ),
    .A2(_04553_),
    .ZN(_04560_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09206_ (.A1(_04448_),
    .A2(_04553_),
    .B(_04560_),
    .ZN(_01227_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09207_ (.A1(\u_cpu.rf_ram.memory[79][7] ),
    .A2(_04553_),
    .ZN(_04561_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09208_ (.A1(_04450_),
    .A2(_04553_),
    .B(_04561_),
    .ZN(_01228_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09209_ (.A1(_02838_),
    .A2(_04349_),
    .ZN(_04562_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09210_ (.I(_04562_),
    .Z(_04563_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09211_ (.A1(\u_cpu.rf_ram.memory[105][0] ),
    .A2(_04563_),
    .ZN(_04564_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09212_ (.A1(_04434_),
    .A2(_04563_),
    .B(_04564_),
    .ZN(_01229_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09213_ (.A1(\u_cpu.rf_ram.memory[105][1] ),
    .A2(_04563_),
    .ZN(_04565_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09214_ (.A1(_04438_),
    .A2(_04563_),
    .B(_04565_),
    .ZN(_01230_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09215_ (.A1(\u_cpu.rf_ram.memory[105][2] ),
    .A2(_04563_),
    .ZN(_04566_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09216_ (.A1(_04440_),
    .A2(_04563_),
    .B(_04566_),
    .ZN(_01231_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09217_ (.A1(\u_cpu.rf_ram.memory[105][3] ),
    .A2(_04563_),
    .ZN(_04567_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09218_ (.A1(_04442_),
    .A2(_04563_),
    .B(_04567_),
    .ZN(_01232_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09219_ (.A1(\u_cpu.rf_ram.memory[105][4] ),
    .A2(_04563_),
    .ZN(_04568_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09220_ (.A1(_04444_),
    .A2(_04563_),
    .B(_04568_),
    .ZN(_01233_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09221_ (.A1(\u_cpu.rf_ram.memory[105][5] ),
    .A2(_04563_),
    .ZN(_04569_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09222_ (.A1(_04446_),
    .A2(_04563_),
    .B(_04569_),
    .ZN(_01234_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09223_ (.A1(\u_cpu.rf_ram.memory[105][6] ),
    .A2(_04563_),
    .ZN(_04570_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09224_ (.A1(_04448_),
    .A2(_04563_),
    .B(_04570_),
    .ZN(_01235_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09225_ (.A1(\u_cpu.rf_ram.memory[105][7] ),
    .A2(_04563_),
    .ZN(_04571_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09226_ (.A1(_04450_),
    .A2(_04563_),
    .B(_04571_),
    .ZN(_01236_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09227_ (.A1(_02780_),
    .A2(_04349_),
    .ZN(_04572_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09228_ (.I(_04572_),
    .Z(_04573_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09229_ (.A1(\u_cpu.rf_ram.memory[106][0] ),
    .A2(_04573_),
    .ZN(_04574_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09230_ (.A1(_04434_),
    .A2(_04573_),
    .B(_04574_),
    .ZN(_01237_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09231_ (.A1(\u_cpu.rf_ram.memory[106][1] ),
    .A2(_04573_),
    .ZN(_04575_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09232_ (.A1(_04438_),
    .A2(_04573_),
    .B(_04575_),
    .ZN(_01238_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09233_ (.A1(\u_cpu.rf_ram.memory[106][2] ),
    .A2(_04573_),
    .ZN(_04576_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09234_ (.A1(_04440_),
    .A2(_04573_),
    .B(_04576_),
    .ZN(_01239_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09235_ (.A1(\u_cpu.rf_ram.memory[106][3] ),
    .A2(_04573_),
    .ZN(_04577_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09236_ (.A1(_04442_),
    .A2(_04573_),
    .B(_04577_),
    .ZN(_01240_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09237_ (.A1(\u_cpu.rf_ram.memory[106][4] ),
    .A2(_04573_),
    .ZN(_04578_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09238_ (.A1(_04444_),
    .A2(_04573_),
    .B(_04578_),
    .ZN(_01241_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09239_ (.A1(\u_cpu.rf_ram.memory[106][5] ),
    .A2(_04573_),
    .ZN(_04579_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09240_ (.A1(_04446_),
    .A2(_04573_),
    .B(_04579_),
    .ZN(_01242_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09241_ (.A1(\u_cpu.rf_ram.memory[106][6] ),
    .A2(_04573_),
    .ZN(_04580_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09242_ (.A1(_04448_),
    .A2(_04573_),
    .B(_04580_),
    .ZN(_01243_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09243_ (.A1(\u_cpu.rf_ram.memory[106][7] ),
    .A2(_04573_),
    .ZN(_04581_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09244_ (.A1(_04450_),
    .A2(_04573_),
    .B(_04581_),
    .ZN(_01244_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09245_ (.A1(_02849_),
    .A2(_04349_),
    .ZN(_04582_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09246_ (.I(_04582_),
    .Z(_04583_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09247_ (.A1(\u_cpu.rf_ram.memory[107][0] ),
    .A2(_04583_),
    .ZN(_04584_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09248_ (.A1(_04434_),
    .A2(_04583_),
    .B(_04584_),
    .ZN(_01245_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09249_ (.A1(\u_cpu.rf_ram.memory[107][1] ),
    .A2(_04583_),
    .ZN(_04585_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09250_ (.A1(_04438_),
    .A2(_04583_),
    .B(_04585_),
    .ZN(_01246_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09251_ (.A1(\u_cpu.rf_ram.memory[107][2] ),
    .A2(_04583_),
    .ZN(_04586_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09252_ (.A1(_04440_),
    .A2(_04583_),
    .B(_04586_),
    .ZN(_01247_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09253_ (.A1(\u_cpu.rf_ram.memory[107][3] ),
    .A2(_04583_),
    .ZN(_04587_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09254_ (.A1(_04442_),
    .A2(_04583_),
    .B(_04587_),
    .ZN(_01248_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09255_ (.A1(\u_cpu.rf_ram.memory[107][4] ),
    .A2(_04583_),
    .ZN(_04588_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09256_ (.A1(_04444_),
    .A2(_04583_),
    .B(_04588_),
    .ZN(_01249_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09257_ (.A1(\u_cpu.rf_ram.memory[107][5] ),
    .A2(_04583_),
    .ZN(_04589_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09258_ (.A1(_04446_),
    .A2(_04583_),
    .B(_04589_),
    .ZN(_01250_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09259_ (.A1(\u_cpu.rf_ram.memory[107][6] ),
    .A2(_04583_),
    .ZN(_04590_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09260_ (.A1(_04448_),
    .A2(_04583_),
    .B(_04590_),
    .ZN(_01251_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09261_ (.A1(\u_cpu.rf_ram.memory[107][7] ),
    .A2(_04583_),
    .ZN(_04591_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09262_ (.A1(_04450_),
    .A2(_04583_),
    .B(_04591_),
    .ZN(_01252_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09263_ (.A1(_02626_),
    .A2(_02825_),
    .ZN(_04592_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09264_ (.I(_04592_),
    .Z(_04593_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09265_ (.A1(\u_cpu.rf_ram.memory[83][0] ),
    .A2(_04593_),
    .ZN(_04594_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09266_ (.A1(_04434_),
    .A2(_04593_),
    .B(_04594_),
    .ZN(_01253_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09267_ (.A1(\u_cpu.rf_ram.memory[83][1] ),
    .A2(_04593_),
    .ZN(_04595_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09268_ (.A1(_04438_),
    .A2(_04593_),
    .B(_04595_),
    .ZN(_01254_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09269_ (.A1(\u_cpu.rf_ram.memory[83][2] ),
    .A2(_04593_),
    .ZN(_04596_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09270_ (.A1(_04440_),
    .A2(_04593_),
    .B(_04596_),
    .ZN(_01255_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09271_ (.A1(\u_cpu.rf_ram.memory[83][3] ),
    .A2(_04593_),
    .ZN(_04597_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09272_ (.A1(_04442_),
    .A2(_04593_),
    .B(_04597_),
    .ZN(_01256_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09273_ (.A1(\u_cpu.rf_ram.memory[83][4] ),
    .A2(_04593_),
    .ZN(_04598_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09274_ (.A1(_04444_),
    .A2(_04593_),
    .B(_04598_),
    .ZN(_01257_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09275_ (.A1(\u_cpu.rf_ram.memory[83][5] ),
    .A2(_04593_),
    .ZN(_04599_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09276_ (.A1(_04446_),
    .A2(_04593_),
    .B(_04599_),
    .ZN(_01258_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09277_ (.A1(\u_cpu.rf_ram.memory[83][6] ),
    .A2(_04593_),
    .ZN(_04600_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09278_ (.A1(_04448_),
    .A2(_04593_),
    .B(_04600_),
    .ZN(_01259_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09279_ (.A1(\u_cpu.rf_ram.memory[83][7] ),
    .A2(_04593_),
    .ZN(_04601_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09280_ (.A1(_04450_),
    .A2(_04593_),
    .B(_04601_),
    .ZN(_01260_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09281_ (.A1(_02814_),
    .A2(_04349_),
    .ZN(_04602_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09282_ (.I(_04602_),
    .Z(_04603_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09283_ (.A1(\u_cpu.rf_ram.memory[108][0] ),
    .A2(_04603_),
    .ZN(_04604_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09284_ (.A1(_04434_),
    .A2(_04603_),
    .B(_04604_),
    .ZN(_01261_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09285_ (.A1(\u_cpu.rf_ram.memory[108][1] ),
    .A2(_04603_),
    .ZN(_04605_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09286_ (.A1(_04438_),
    .A2(_04603_),
    .B(_04605_),
    .ZN(_01262_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09287_ (.A1(\u_cpu.rf_ram.memory[108][2] ),
    .A2(_04603_),
    .ZN(_04606_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09288_ (.A1(_04440_),
    .A2(_04603_),
    .B(_04606_),
    .ZN(_01263_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09289_ (.A1(\u_cpu.rf_ram.memory[108][3] ),
    .A2(_04603_),
    .ZN(_04607_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09290_ (.A1(_04442_),
    .A2(_04603_),
    .B(_04607_),
    .ZN(_01264_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09291_ (.A1(\u_cpu.rf_ram.memory[108][4] ),
    .A2(_04603_),
    .ZN(_04608_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09292_ (.A1(_04444_),
    .A2(_04603_),
    .B(_04608_),
    .ZN(_01265_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09293_ (.A1(\u_cpu.rf_ram.memory[108][5] ),
    .A2(_04603_),
    .ZN(_04609_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09294_ (.A1(_04446_),
    .A2(_04603_),
    .B(_04609_),
    .ZN(_01266_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09295_ (.A1(\u_cpu.rf_ram.memory[108][6] ),
    .A2(_04603_),
    .ZN(_04610_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09296_ (.A1(_04448_),
    .A2(_04603_),
    .B(_04610_),
    .ZN(_01267_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09297_ (.A1(\u_cpu.rf_ram.memory[108][7] ),
    .A2(_04603_),
    .ZN(_04611_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09298_ (.A1(_04450_),
    .A2(_04603_),
    .B(_04611_),
    .ZN(_01268_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09299_ (.A1(_02675_),
    .A2(_02768_),
    .ZN(_04612_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09300_ (.I(_04612_),
    .Z(_04613_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09301_ (.A1(\u_cpu.rf_ram.memory[69][0] ),
    .A2(_04613_),
    .ZN(_04614_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09302_ (.A1(_04434_),
    .A2(_04613_),
    .B(_04614_),
    .ZN(_01269_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09303_ (.A1(\u_cpu.rf_ram.memory[69][1] ),
    .A2(_04613_),
    .ZN(_04615_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09304_ (.A1(_04438_),
    .A2(_04613_),
    .B(_04615_),
    .ZN(_01270_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09305_ (.A1(\u_cpu.rf_ram.memory[69][2] ),
    .A2(_04613_),
    .ZN(_04616_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09306_ (.A1(_04440_),
    .A2(_04613_),
    .B(_04616_),
    .ZN(_01271_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09307_ (.A1(\u_cpu.rf_ram.memory[69][3] ),
    .A2(_04613_),
    .ZN(_04617_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09308_ (.A1(_04442_),
    .A2(_04613_),
    .B(_04617_),
    .ZN(_01272_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09309_ (.A1(\u_cpu.rf_ram.memory[69][4] ),
    .A2(_04613_),
    .ZN(_04618_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09310_ (.A1(_04444_),
    .A2(_04613_),
    .B(_04618_),
    .ZN(_01273_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09311_ (.A1(\u_cpu.rf_ram.memory[69][5] ),
    .A2(_04613_),
    .ZN(_04619_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09312_ (.A1(_04446_),
    .A2(_04613_),
    .B(_04619_),
    .ZN(_01274_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09313_ (.A1(\u_cpu.rf_ram.memory[69][6] ),
    .A2(_04613_),
    .ZN(_04620_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09314_ (.A1(_04448_),
    .A2(_04613_),
    .B(_04620_),
    .ZN(_01275_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09315_ (.A1(\u_cpu.rf_ram.memory[69][7] ),
    .A2(_04613_),
    .ZN(_04621_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09316_ (.A1(_04450_),
    .A2(_04613_),
    .B(_04621_),
    .ZN(_01276_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09317_ (.I(_02631_),
    .Z(_04622_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09318_ (.A1(_02626_),
    .A2(_02717_),
    .ZN(_04623_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09319_ (.I(_04623_),
    .Z(_04624_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09320_ (.A1(\u_cpu.rf_ram.memory[84][0] ),
    .A2(_04624_),
    .ZN(_04625_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09321_ (.A1(_04622_),
    .A2(_04624_),
    .B(_04625_),
    .ZN(_01277_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09322_ (.I(_02636_),
    .Z(_04626_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09323_ (.A1(\u_cpu.rf_ram.memory[84][1] ),
    .A2(_04624_),
    .ZN(_04627_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09324_ (.A1(_04626_),
    .A2(_04624_),
    .B(_04627_),
    .ZN(_01278_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09325_ (.I(_02641_),
    .Z(_04628_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09326_ (.A1(\u_cpu.rf_ram.memory[84][2] ),
    .A2(_04624_),
    .ZN(_04629_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09327_ (.A1(_04628_),
    .A2(_04624_),
    .B(_04629_),
    .ZN(_01279_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09328_ (.I(_02646_),
    .Z(_04630_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09329_ (.A1(\u_cpu.rf_ram.memory[84][3] ),
    .A2(_04624_),
    .ZN(_04631_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09330_ (.A1(_04630_),
    .A2(_04624_),
    .B(_04631_),
    .ZN(_01280_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09331_ (.I(_02651_),
    .Z(_04632_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09332_ (.A1(\u_cpu.rf_ram.memory[84][4] ),
    .A2(_04624_),
    .ZN(_04633_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09333_ (.A1(_04632_),
    .A2(_04624_),
    .B(_04633_),
    .ZN(_01281_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09334_ (.I(_02656_),
    .Z(_04634_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09335_ (.A1(\u_cpu.rf_ram.memory[84][5] ),
    .A2(_04624_),
    .ZN(_04635_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09336_ (.A1(_04634_),
    .A2(_04624_),
    .B(_04635_),
    .ZN(_01282_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09337_ (.I(_02661_),
    .Z(_04636_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09338_ (.A1(\u_cpu.rf_ram.memory[84][6] ),
    .A2(_04624_),
    .ZN(_04637_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09339_ (.A1(_04636_),
    .A2(_04624_),
    .B(_04637_),
    .ZN(_01283_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09340_ (.I(_02666_),
    .Z(_04638_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09341_ (.A1(\u_cpu.rf_ram.memory[84][7] ),
    .A2(_04624_),
    .ZN(_04639_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09342_ (.A1(_04638_),
    .A2(_04624_),
    .B(_04639_),
    .ZN(_01284_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09343_ (.A1(_02827_),
    .A2(_02849_),
    .ZN(_04640_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09344_ (.I(_04640_),
    .Z(_04641_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09345_ (.A1(\u_cpu.rf_ram.memory[59][0] ),
    .A2(_04641_),
    .ZN(_04642_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09346_ (.A1(_04622_),
    .A2(_04641_),
    .B(_04642_),
    .ZN(_01285_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09347_ (.A1(\u_cpu.rf_ram.memory[59][1] ),
    .A2(_04641_),
    .ZN(_04643_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09348_ (.A1(_04626_),
    .A2(_04641_),
    .B(_04643_),
    .ZN(_01286_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09349_ (.A1(\u_cpu.rf_ram.memory[59][2] ),
    .A2(_04641_),
    .ZN(_04644_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09350_ (.A1(_04628_),
    .A2(_04641_),
    .B(_04644_),
    .ZN(_01287_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09351_ (.A1(\u_cpu.rf_ram.memory[59][3] ),
    .A2(_04641_),
    .ZN(_04645_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09352_ (.A1(_04630_),
    .A2(_04641_),
    .B(_04645_),
    .ZN(_01288_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09353_ (.A1(\u_cpu.rf_ram.memory[59][4] ),
    .A2(_04641_),
    .ZN(_04646_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09354_ (.A1(_04632_),
    .A2(_04641_),
    .B(_04646_),
    .ZN(_01289_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09355_ (.A1(\u_cpu.rf_ram.memory[59][5] ),
    .A2(_04641_),
    .ZN(_04647_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09356_ (.A1(_04634_),
    .A2(_04641_),
    .B(_04647_),
    .ZN(_01290_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09357_ (.A1(\u_cpu.rf_ram.memory[59][6] ),
    .A2(_04641_),
    .ZN(_04648_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09358_ (.A1(_04636_),
    .A2(_04641_),
    .B(_04648_),
    .ZN(_01291_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09359_ (.A1(\u_cpu.rf_ram.memory[59][7] ),
    .A2(_04641_),
    .ZN(_04649_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09360_ (.A1(_04638_),
    .A2(_04641_),
    .B(_04649_),
    .ZN(_01292_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09361_ (.A1(_02731_),
    .A2(_02780_),
    .ZN(_04650_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09362_ (.I(_04650_),
    .ZN(_04651_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09363_ (.A1(\u_cpu.rf_ram.memory[10][0] ),
    .A2(_04651_),
    .ZN(_04652_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09364_ (.A1(_02632_),
    .A2(_04651_),
    .B(_04652_),
    .ZN(_01293_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09365_ (.A1(\u_cpu.rf_ram.memory[10][1] ),
    .A2(_04651_),
    .ZN(_04653_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09366_ (.A1(_02637_),
    .A2(_04651_),
    .B(_04653_),
    .ZN(_01294_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09367_ (.A1(\u_cpu.rf_ram.memory[10][2] ),
    .A2(_04651_),
    .ZN(_04654_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09368_ (.A1(_02642_),
    .A2(_04651_),
    .B(_04654_),
    .ZN(_01295_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09369_ (.A1(\u_cpu.rf_ram.memory[10][3] ),
    .A2(_04651_),
    .ZN(_04655_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09370_ (.A1(_02647_),
    .A2(_04651_),
    .B(_04655_),
    .ZN(_01296_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09371_ (.A1(\u_cpu.rf_ram.memory[10][4] ),
    .A2(_04651_),
    .ZN(_04656_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09372_ (.A1(_02652_),
    .A2(_04651_),
    .B(_04656_),
    .ZN(_01297_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09373_ (.A1(\u_cpu.rf_ram.memory[10][5] ),
    .A2(_04651_),
    .ZN(_04657_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09374_ (.A1(_02657_),
    .A2(_04651_),
    .B(_04657_),
    .ZN(_01298_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09375_ (.A1(\u_cpu.rf_ram.memory[10][6] ),
    .A2(_04651_),
    .ZN(_04658_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09376_ (.A1(_02662_),
    .A2(_04651_),
    .B(_04658_),
    .ZN(_01299_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09377_ (.A1(\u_cpu.rf_ram.memory[10][7] ),
    .A2(_04651_),
    .ZN(_04659_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09378_ (.A1(_02667_),
    .A2(_04651_),
    .B(_04659_),
    .ZN(_01300_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09379_ (.A1(_02626_),
    .A2(_02675_),
    .ZN(_04660_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09380_ (.I(_04660_),
    .Z(_04661_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09381_ (.A1(\u_cpu.rf_ram.memory[85][0] ),
    .A2(_04661_),
    .ZN(_04662_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09382_ (.A1(_04622_),
    .A2(_04661_),
    .B(_04662_),
    .ZN(_01301_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09383_ (.A1(\u_cpu.rf_ram.memory[85][1] ),
    .A2(_04661_),
    .ZN(_04663_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09384_ (.A1(_04626_),
    .A2(_04661_),
    .B(_04663_),
    .ZN(_01302_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09385_ (.A1(\u_cpu.rf_ram.memory[85][2] ),
    .A2(_04661_),
    .ZN(_04664_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09386_ (.A1(_04628_),
    .A2(_04661_),
    .B(_04664_),
    .ZN(_01303_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09387_ (.A1(\u_cpu.rf_ram.memory[85][3] ),
    .A2(_04661_),
    .ZN(_04665_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09388_ (.A1(_04630_),
    .A2(_04661_),
    .B(_04665_),
    .ZN(_01304_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09389_ (.A1(\u_cpu.rf_ram.memory[85][4] ),
    .A2(_04661_),
    .ZN(_04666_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09390_ (.A1(_04632_),
    .A2(_04661_),
    .B(_04666_),
    .ZN(_01305_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09391_ (.A1(\u_cpu.rf_ram.memory[85][5] ),
    .A2(_04661_),
    .ZN(_04667_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09392_ (.A1(_04634_),
    .A2(_04661_),
    .B(_04667_),
    .ZN(_01306_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09393_ (.A1(\u_cpu.rf_ram.memory[85][6] ),
    .A2(_04661_),
    .ZN(_04668_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09394_ (.A1(_04636_),
    .A2(_04661_),
    .B(_04668_),
    .ZN(_01307_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09395_ (.A1(\u_cpu.rf_ram.memory[85][7] ),
    .A2(_04661_),
    .ZN(_04669_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09396_ (.A1(_04638_),
    .A2(_04661_),
    .B(_04669_),
    .ZN(_01308_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09397_ (.A1(_02766_),
    .A2(_04349_),
    .ZN(_04670_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09398_ (.I(_04670_),
    .Z(_04671_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09399_ (.A1(\u_cpu.rf_ram.memory[110][0] ),
    .A2(_04671_),
    .ZN(_04672_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09400_ (.A1(_04622_),
    .A2(_04671_),
    .B(_04672_),
    .ZN(_01309_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09401_ (.A1(\u_cpu.rf_ram.memory[110][1] ),
    .A2(_04671_),
    .ZN(_04673_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09402_ (.A1(_04626_),
    .A2(_04671_),
    .B(_04673_),
    .ZN(_01310_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09403_ (.A1(\u_cpu.rf_ram.memory[110][2] ),
    .A2(_04671_),
    .ZN(_04674_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09404_ (.A1(_04628_),
    .A2(_04671_),
    .B(_04674_),
    .ZN(_01311_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09405_ (.A1(\u_cpu.rf_ram.memory[110][3] ),
    .A2(_04671_),
    .ZN(_04675_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09406_ (.A1(_04630_),
    .A2(_04671_),
    .B(_04675_),
    .ZN(_01312_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09407_ (.A1(\u_cpu.rf_ram.memory[110][4] ),
    .A2(_04671_),
    .ZN(_04676_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09408_ (.A1(_04632_),
    .A2(_04671_),
    .B(_04676_),
    .ZN(_01313_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09409_ (.A1(\u_cpu.rf_ram.memory[110][5] ),
    .A2(_04671_),
    .ZN(_04677_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09410_ (.A1(_04634_),
    .A2(_04671_),
    .B(_04677_),
    .ZN(_01314_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09411_ (.A1(\u_cpu.rf_ram.memory[110][6] ),
    .A2(_04671_),
    .ZN(_04678_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09412_ (.A1(_04636_),
    .A2(_04671_),
    .B(_04678_),
    .ZN(_01315_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09413_ (.A1(\u_cpu.rf_ram.memory[110][7] ),
    .A2(_04671_),
    .ZN(_04679_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09414_ (.A1(_04638_),
    .A2(_04671_),
    .B(_04679_),
    .ZN(_01316_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09415_ (.A1(_02626_),
    .A2(_03037_),
    .ZN(_04680_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09416_ (.I(_04680_),
    .Z(_04681_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09417_ (.A1(\u_cpu.rf_ram.memory[86][0] ),
    .A2(_04681_),
    .ZN(_04682_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09418_ (.A1(_04622_),
    .A2(_04681_),
    .B(_04682_),
    .ZN(_01317_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09419_ (.A1(\u_cpu.rf_ram.memory[86][1] ),
    .A2(_04681_),
    .ZN(_04683_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09420_ (.A1(_04626_),
    .A2(_04681_),
    .B(_04683_),
    .ZN(_01318_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09421_ (.A1(\u_cpu.rf_ram.memory[86][2] ),
    .A2(_04681_),
    .ZN(_04684_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09422_ (.A1(_04628_),
    .A2(_04681_),
    .B(_04684_),
    .ZN(_01319_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09423_ (.A1(\u_cpu.rf_ram.memory[86][3] ),
    .A2(_04681_),
    .ZN(_04685_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09424_ (.A1(_04630_),
    .A2(_04681_),
    .B(_04685_),
    .ZN(_01320_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09425_ (.A1(\u_cpu.rf_ram.memory[86][4] ),
    .A2(_04681_),
    .ZN(_04686_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09426_ (.A1(_04632_),
    .A2(_04681_),
    .B(_04686_),
    .ZN(_01321_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09427_ (.A1(\u_cpu.rf_ram.memory[86][5] ),
    .A2(_04681_),
    .ZN(_04687_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09428_ (.A1(_04634_),
    .A2(_04681_),
    .B(_04687_),
    .ZN(_01322_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09429_ (.A1(\u_cpu.rf_ram.memory[86][6] ),
    .A2(_04681_),
    .ZN(_04688_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09430_ (.A1(_04636_),
    .A2(_04681_),
    .B(_04688_),
    .ZN(_01323_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09431_ (.A1(\u_cpu.rf_ram.memory[86][7] ),
    .A2(_04681_),
    .ZN(_04689_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09432_ (.A1(_04638_),
    .A2(_04681_),
    .B(_04689_),
    .ZN(_01324_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09433_ (.A1(_02870_),
    .A2(_04349_),
    .ZN(_04690_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09434_ (.I(_04690_),
    .Z(_04691_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09435_ (.A1(\u_cpu.rf_ram.memory[111][0] ),
    .A2(_04691_),
    .ZN(_04692_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09436_ (.A1(_04622_),
    .A2(_04691_),
    .B(_04692_),
    .ZN(_01325_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09437_ (.A1(\u_cpu.rf_ram.memory[111][1] ),
    .A2(_04691_),
    .ZN(_04693_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09438_ (.A1(_04626_),
    .A2(_04691_),
    .B(_04693_),
    .ZN(_01326_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09439_ (.A1(\u_cpu.rf_ram.memory[111][2] ),
    .A2(_04691_),
    .ZN(_04694_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09440_ (.A1(_04628_),
    .A2(_04691_),
    .B(_04694_),
    .ZN(_01327_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09441_ (.A1(\u_cpu.rf_ram.memory[111][3] ),
    .A2(_04691_),
    .ZN(_04695_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09442_ (.A1(_04630_),
    .A2(_04691_),
    .B(_04695_),
    .ZN(_01328_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09443_ (.A1(\u_cpu.rf_ram.memory[111][4] ),
    .A2(_04691_),
    .ZN(_04696_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09444_ (.A1(_04632_),
    .A2(_04691_),
    .B(_04696_),
    .ZN(_01329_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09445_ (.A1(\u_cpu.rf_ram.memory[111][5] ),
    .A2(_04691_),
    .ZN(_04697_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09446_ (.A1(_04634_),
    .A2(_04691_),
    .B(_04697_),
    .ZN(_01330_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09447_ (.A1(\u_cpu.rf_ram.memory[111][6] ),
    .A2(_04691_),
    .ZN(_04698_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09448_ (.A1(_04636_),
    .A2(_04691_),
    .B(_04698_),
    .ZN(_01331_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09449_ (.A1(\u_cpu.rf_ram.memory[111][7] ),
    .A2(_04691_),
    .ZN(_04699_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09450_ (.A1(_04638_),
    .A2(_04691_),
    .B(_04699_),
    .ZN(_01332_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09451_ (.A1(_02626_),
    .A2(_02743_),
    .ZN(_04700_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09452_ (.I(_04700_),
    .Z(_04701_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09453_ (.A1(\u_cpu.rf_ram.memory[87][0] ),
    .A2(_04701_),
    .ZN(_04702_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09454_ (.A1(_04622_),
    .A2(_04701_),
    .B(_04702_),
    .ZN(_01333_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09455_ (.A1(\u_cpu.rf_ram.memory[87][1] ),
    .A2(_04701_),
    .ZN(_04703_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09456_ (.A1(_04626_),
    .A2(_04701_),
    .B(_04703_),
    .ZN(_01334_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09457_ (.A1(\u_cpu.rf_ram.memory[87][2] ),
    .A2(_04701_),
    .ZN(_04704_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09458_ (.A1(_04628_),
    .A2(_04701_),
    .B(_04704_),
    .ZN(_01335_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09459_ (.A1(\u_cpu.rf_ram.memory[87][3] ),
    .A2(_04701_),
    .ZN(_04705_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09460_ (.A1(_04630_),
    .A2(_04701_),
    .B(_04705_),
    .ZN(_01336_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09461_ (.A1(\u_cpu.rf_ram.memory[87][4] ),
    .A2(_04701_),
    .ZN(_04706_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09462_ (.A1(_04632_),
    .A2(_04701_),
    .B(_04706_),
    .ZN(_01337_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09463_ (.A1(\u_cpu.rf_ram.memory[87][5] ),
    .A2(_04701_),
    .ZN(_04707_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09464_ (.A1(_04634_),
    .A2(_04701_),
    .B(_04707_),
    .ZN(_01338_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09465_ (.A1(\u_cpu.rf_ram.memory[87][6] ),
    .A2(_04701_),
    .ZN(_04708_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09466_ (.A1(_04636_),
    .A2(_04701_),
    .B(_04708_),
    .ZN(_01339_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09467_ (.A1(\u_cpu.rf_ram.memory[87][7] ),
    .A2(_04701_),
    .ZN(_04709_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09468_ (.A1(_04638_),
    .A2(_04701_),
    .B(_04709_),
    .ZN(_01340_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09469_ (.A1(_02626_),
    .A2(_02954_),
    .ZN(_04710_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09470_ (.I(_04710_),
    .Z(_04711_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09471_ (.A1(\u_cpu.rf_ram.memory[88][0] ),
    .A2(_04711_),
    .ZN(_04712_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09472_ (.A1(_04622_),
    .A2(_04711_),
    .B(_04712_),
    .ZN(_01341_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09473_ (.A1(\u_cpu.rf_ram.memory[88][1] ),
    .A2(_04711_),
    .ZN(_04713_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09474_ (.A1(_04626_),
    .A2(_04711_),
    .B(_04713_),
    .ZN(_01342_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09475_ (.A1(\u_cpu.rf_ram.memory[88][2] ),
    .A2(_04711_),
    .ZN(_04714_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09476_ (.A1(_04628_),
    .A2(_04711_),
    .B(_04714_),
    .ZN(_01343_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09477_ (.A1(\u_cpu.rf_ram.memory[88][3] ),
    .A2(_04711_),
    .ZN(_04715_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09478_ (.A1(_04630_),
    .A2(_04711_),
    .B(_04715_),
    .ZN(_01344_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09479_ (.A1(\u_cpu.rf_ram.memory[88][4] ),
    .A2(_04711_),
    .ZN(_04716_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09480_ (.A1(_04632_),
    .A2(_04711_),
    .B(_04716_),
    .ZN(_01345_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09481_ (.A1(\u_cpu.rf_ram.memory[88][5] ),
    .A2(_04711_),
    .ZN(_04717_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09482_ (.A1(_04634_),
    .A2(_04711_),
    .B(_04717_),
    .ZN(_01346_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09483_ (.A1(\u_cpu.rf_ram.memory[88][6] ),
    .A2(_04711_),
    .ZN(_04718_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09484_ (.A1(_04636_),
    .A2(_04711_),
    .B(_04718_),
    .ZN(_01347_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09485_ (.A1(\u_cpu.rf_ram.memory[88][7] ),
    .A2(_04711_),
    .ZN(_04719_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09486_ (.A1(_04638_),
    .A2(_04711_),
    .B(_04719_),
    .ZN(_01348_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09487_ (.A1(_02263_),
    .A2(_02303_),
    .ZN(_04720_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09488_ (.A1(_02259_),
    .A2(_02297_),
    .A3(_02292_),
    .ZN(_04721_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09489_ (.A1(_04720_),
    .A2(_04721_),
    .Z(_04722_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09490_ (.I(_04722_),
    .Z(_04723_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09491_ (.I(\u_cpu.cpu.genblk3.csr.mcause3_0[1] ),
    .ZN(_04724_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _09492_ (.A1(\u_cpu.cpu.decode.op21 ),
    .A2(_01443_),
    .A3(_01457_),
    .ZN(_04725_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09493_ (.A1(\u_cpu.cpu.genblk3.csr.o_new_irq ),
    .A2(_04725_),
    .ZN(_04726_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09494_ (.A1(\u_cpu.cpu.state.genblk1.misalign_trap_sync_r ),
    .A2(_04724_),
    .B(_04726_),
    .ZN(_04727_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09495_ (.A1(_04723_),
    .A2(_04727_),
    .ZN(_04728_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09496_ (.A1(_02295_),
    .A2(_04723_),
    .B(_04728_),
    .ZN(_01349_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09497_ (.I(\u_cpu.cpu.genblk3.csr.mcause3_0[2] ),
    .ZN(_04729_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _09498_ (.A1(_02305_),
    .A2(_02400_),
    .B1(_04729_),
    .B2(\u_cpu.cpu.state.genblk1.misalign_trap_sync_r ),
    .C(_04726_),
    .ZN(_04730_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09499_ (.A1(_04723_),
    .A2(_04730_),
    .ZN(_04731_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09500_ (.A1(_04724_),
    .A2(_04723_),
    .B(_04731_),
    .ZN(_01350_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09501_ (.I(\u_cpu.cpu.genblk3.csr.mcause3_0[3] ),
    .ZN(_04732_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09502_ (.A1(_04732_),
    .A2(_02303_),
    .B(_01458_),
    .C(_02305_),
    .ZN(_04733_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09503_ (.I0(_04733_),
    .I1(\u_cpu.cpu.genblk3.csr.mcause3_0[2] ),
    .S(_04723_),
    .Z(_04734_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09504_ (.I(_04734_),
    .Z(_01351_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09505_ (.A1(_02325_),
    .A2(_04725_),
    .B(_04723_),
    .ZN(_04735_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09506_ (.A1(_04732_),
    .A2(_04723_),
    .B1(_04735_),
    .B2(_02302_),
    .ZN(_01352_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09507_ (.A1(_01458_),
    .A2(_02302_),
    .ZN(_04736_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09508_ (.A1(_02263_),
    .A2(_02297_),
    .B(_02303_),
    .ZN(_04737_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09509_ (.I0(_04736_),
    .I1(\u_cpu.cpu.genblk3.csr.mcause31 ),
    .S(_04737_),
    .Z(_04738_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09510_ (.I(_04738_),
    .Z(_01353_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09511_ (.I(\u_cpu.cpu.genblk3.csr.mstatus_mpie ),
    .ZN(_04739_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09512_ (.A1(\u_cpu.cpu.genblk3.csr.mstatus_mie ),
    .A2(_04720_),
    .ZN(_04740_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09513_ (.A1(_04739_),
    .A2(_04720_),
    .B(_04740_),
    .ZN(_01354_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09514_ (.I(\u_cpu.cpu.genblk3.csr.mie_mtie ),
    .ZN(_04741_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _09515_ (.A1(\u_cpu.cpu.decode.co_ebreak ),
    .A2(\u_cpu.cpu.mem_bytecnt[1] ),
    .A3(_02291_),
    .A4(_02290_),
    .ZN(_04742_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09516_ (.A1(_02293_),
    .A2(_03605_),
    .A3(_04742_),
    .ZN(_04743_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09517_ (.A1(_02301_),
    .A2(_04743_),
    .B(_02396_),
    .ZN(_04744_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09518_ (.A1(_04741_),
    .A2(_04743_),
    .B(_04744_),
    .ZN(_01355_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09519_ (.A1(_01477_),
    .A2(_02294_),
    .ZN(_04745_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09520_ (.A1(_04739_),
    .A2(_01477_),
    .B(_02303_),
    .C(_04745_),
    .ZN(_04746_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09521_ (.A1(_01477_),
    .A2(_02301_),
    .B(_04746_),
    .ZN(_04747_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09522_ (.A1(\u_cpu.cpu.genblk3.csr.mstatus_mie ),
    .A2(_04720_),
    .A3(_04745_),
    .ZN(_04748_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09523_ (.A1(_04747_),
    .A2(_04748_),
    .ZN(_01356_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09524_ (.A1(\u_cpu.cpu.ctrl.i_iscomp ),
    .A2(_03897_),
    .ZN(_04749_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09525_ (.A1(_03966_),
    .A2(_04749_),
    .ZN(_01357_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09526_ (.A1(\u_cpu.cpu.genblk3.csr.o_new_irq ),
    .A2(_03611_),
    .ZN(_04750_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _09527_ (.A1(_02395_),
    .A2(\u_cpu.cpu.genblk3.csr.timer_irq_r ),
    .A3(_04235_),
    .B(_04750_),
    .ZN(_01358_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09528_ (.A1(_02677_),
    .A2(_02849_),
    .ZN(_04751_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09529_ (.I(_04751_),
    .Z(_04752_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09530_ (.A1(\u_cpu.rf_ram.memory[27][0] ),
    .A2(_04752_),
    .ZN(_04753_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09531_ (.A1(_04622_),
    .A2(_04752_),
    .B(_04753_),
    .ZN(_01359_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09532_ (.A1(\u_cpu.rf_ram.memory[27][1] ),
    .A2(_04752_),
    .ZN(_04754_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09533_ (.A1(_04626_),
    .A2(_04752_),
    .B(_04754_),
    .ZN(_01360_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09534_ (.A1(\u_cpu.rf_ram.memory[27][2] ),
    .A2(_04752_),
    .ZN(_04755_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09535_ (.A1(_04628_),
    .A2(_04752_),
    .B(_04755_),
    .ZN(_01361_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09536_ (.A1(\u_cpu.rf_ram.memory[27][3] ),
    .A2(_04752_),
    .ZN(_04756_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09537_ (.A1(_04630_),
    .A2(_04752_),
    .B(_04756_),
    .ZN(_01362_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09538_ (.A1(\u_cpu.rf_ram.memory[27][4] ),
    .A2(_04752_),
    .ZN(_04757_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09539_ (.A1(_04632_),
    .A2(_04752_),
    .B(_04757_),
    .ZN(_01363_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09540_ (.A1(\u_cpu.rf_ram.memory[27][5] ),
    .A2(_04752_),
    .ZN(_04758_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09541_ (.A1(_04634_),
    .A2(_04752_),
    .B(_04758_),
    .ZN(_01364_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09542_ (.A1(\u_cpu.rf_ram.memory[27][6] ),
    .A2(_04752_),
    .ZN(_04759_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09543_ (.A1(_04636_),
    .A2(_04752_),
    .B(_04759_),
    .ZN(_01365_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09544_ (.A1(\u_cpu.rf_ram.memory[27][7] ),
    .A2(_04752_),
    .ZN(_04760_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09545_ (.A1(_04638_),
    .A2(_04752_),
    .B(_04760_),
    .ZN(_01366_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09546_ (.A1(_02677_),
    .A2(_02780_),
    .ZN(_04761_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09547_ (.I(_04761_),
    .Z(_04762_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09548_ (.A1(\u_cpu.rf_ram.memory[26][0] ),
    .A2(_04762_),
    .ZN(_04763_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09549_ (.A1(_04622_),
    .A2(_04762_),
    .B(_04763_),
    .ZN(_01367_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09550_ (.A1(\u_cpu.rf_ram.memory[26][1] ),
    .A2(_04762_),
    .ZN(_04764_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09551_ (.A1(_04626_),
    .A2(_04762_),
    .B(_04764_),
    .ZN(_01368_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09552_ (.A1(\u_cpu.rf_ram.memory[26][2] ),
    .A2(_04762_),
    .ZN(_04765_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09553_ (.A1(_04628_),
    .A2(_04762_),
    .B(_04765_),
    .ZN(_01369_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09554_ (.A1(\u_cpu.rf_ram.memory[26][3] ),
    .A2(_04762_),
    .ZN(_04766_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09555_ (.A1(_04630_),
    .A2(_04762_),
    .B(_04766_),
    .ZN(_01370_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09556_ (.A1(\u_cpu.rf_ram.memory[26][4] ),
    .A2(_04762_),
    .ZN(_04767_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09557_ (.A1(_04632_),
    .A2(_04762_),
    .B(_04767_),
    .ZN(_01371_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09558_ (.A1(\u_cpu.rf_ram.memory[26][5] ),
    .A2(_04762_),
    .ZN(_04768_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09559_ (.A1(_04634_),
    .A2(_04762_),
    .B(_04768_),
    .ZN(_01372_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09560_ (.A1(\u_cpu.rf_ram.memory[26][6] ),
    .A2(_04762_),
    .ZN(_04769_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09561_ (.A1(_04636_),
    .A2(_04762_),
    .B(_04769_),
    .ZN(_01373_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09562_ (.A1(\u_cpu.rf_ram.memory[26][7] ),
    .A2(_04762_),
    .ZN(_04770_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09563_ (.A1(_04638_),
    .A2(_04762_),
    .B(_04770_),
    .ZN(_01374_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09564_ (.A1(_02677_),
    .A2(_02838_),
    .ZN(_04771_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09565_ (.I(_04771_),
    .Z(_04772_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09566_ (.A1(\u_cpu.rf_ram.memory[25][0] ),
    .A2(_04772_),
    .ZN(_04773_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09567_ (.A1(_04622_),
    .A2(_04772_),
    .B(_04773_),
    .ZN(_01375_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09568_ (.A1(\u_cpu.rf_ram.memory[25][1] ),
    .A2(_04772_),
    .ZN(_04774_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09569_ (.A1(_04626_),
    .A2(_04772_),
    .B(_04774_),
    .ZN(_01376_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09570_ (.A1(\u_cpu.rf_ram.memory[25][2] ),
    .A2(_04772_),
    .ZN(_04775_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09571_ (.A1(_04628_),
    .A2(_04772_),
    .B(_04775_),
    .ZN(_01377_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09572_ (.A1(\u_cpu.rf_ram.memory[25][3] ),
    .A2(_04772_),
    .ZN(_04776_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09573_ (.A1(_04630_),
    .A2(_04772_),
    .B(_04776_),
    .ZN(_01378_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09574_ (.A1(\u_cpu.rf_ram.memory[25][4] ),
    .A2(_04772_),
    .ZN(_04777_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09575_ (.A1(_04632_),
    .A2(_04772_),
    .B(_04777_),
    .ZN(_01379_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09576_ (.A1(\u_cpu.rf_ram.memory[25][5] ),
    .A2(_04772_),
    .ZN(_04778_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09577_ (.A1(_04634_),
    .A2(_04772_),
    .B(_04778_),
    .ZN(_01380_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09578_ (.A1(\u_cpu.rf_ram.memory[25][6] ),
    .A2(_04772_),
    .ZN(_04779_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09579_ (.A1(_04636_),
    .A2(_04772_),
    .B(_04779_),
    .ZN(_01381_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09580_ (.A1(\u_cpu.rf_ram.memory[25][7] ),
    .A2(_04772_),
    .ZN(_04780_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09581_ (.A1(_04638_),
    .A2(_04772_),
    .B(_04780_),
    .ZN(_01382_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09582_ (.A1(_02677_),
    .A2(_02954_),
    .ZN(_04781_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09583_ (.I(_04781_),
    .Z(_04782_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09584_ (.A1(\u_cpu.rf_ram.memory[24][0] ),
    .A2(_04782_),
    .ZN(_04783_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09585_ (.A1(_04622_),
    .A2(_04782_),
    .B(_04783_),
    .ZN(_01383_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09586_ (.A1(\u_cpu.rf_ram.memory[24][1] ),
    .A2(_04782_),
    .ZN(_04784_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09587_ (.A1(_04626_),
    .A2(_04782_),
    .B(_04784_),
    .ZN(_01384_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09588_ (.A1(\u_cpu.rf_ram.memory[24][2] ),
    .A2(_04782_),
    .ZN(_04785_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09589_ (.A1(_04628_),
    .A2(_04782_),
    .B(_04785_),
    .ZN(_01385_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09590_ (.A1(\u_cpu.rf_ram.memory[24][3] ),
    .A2(_04782_),
    .ZN(_04786_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09591_ (.A1(_04630_),
    .A2(_04782_),
    .B(_04786_),
    .ZN(_01386_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09592_ (.A1(\u_cpu.rf_ram.memory[24][4] ),
    .A2(_04782_),
    .ZN(_04787_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09593_ (.A1(_04632_),
    .A2(_04782_),
    .B(_04787_),
    .ZN(_01387_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09594_ (.A1(\u_cpu.rf_ram.memory[24][5] ),
    .A2(_04782_),
    .ZN(_04788_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09595_ (.A1(_04634_),
    .A2(_04782_),
    .B(_04788_),
    .ZN(_01388_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09596_ (.A1(\u_cpu.rf_ram.memory[24][6] ),
    .A2(_04782_),
    .ZN(_04789_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09597_ (.A1(_04636_),
    .A2(_04782_),
    .B(_04789_),
    .ZN(_01389_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09598_ (.A1(\u_cpu.rf_ram.memory[24][7] ),
    .A2(_04782_),
    .ZN(_04790_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09599_ (.A1(_04638_),
    .A2(_04782_),
    .B(_04790_),
    .ZN(_01390_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09600_ (.A1(_02731_),
    .A2(_02754_),
    .Z(_04791_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09601_ (.I(_04791_),
    .Z(_04792_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09602_ (.A1(\u_cpu.rf_ram.memory[0][0] ),
    .A2(_04792_),
    .ZN(_04793_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09603_ (.A1(_02669_),
    .A2(_04792_),
    .B(_04793_),
    .ZN(_01391_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09604_ (.A1(\u_cpu.rf_ram.memory[0][1] ),
    .A2(_04792_),
    .ZN(_04794_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09605_ (.A1(_02681_),
    .A2(_04792_),
    .B(_04794_),
    .ZN(_01392_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09606_ (.A1(\u_cpu.rf_ram.memory[0][2] ),
    .A2(_04792_),
    .ZN(_04795_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09607_ (.A1(_02683_),
    .A2(_04792_),
    .B(_04795_),
    .ZN(_01393_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09608_ (.A1(\u_cpu.rf_ram.memory[0][3] ),
    .A2(_04792_),
    .ZN(_04796_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09609_ (.A1(_02685_),
    .A2(_04792_),
    .B(_04796_),
    .ZN(_01394_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09610_ (.A1(\u_cpu.rf_ram.memory[0][4] ),
    .A2(_04792_),
    .ZN(_04797_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09611_ (.A1(_02687_),
    .A2(_04792_),
    .B(_04797_),
    .ZN(_01395_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09612_ (.A1(\u_cpu.rf_ram.memory[0][5] ),
    .A2(_04792_),
    .ZN(_04798_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09613_ (.A1(_02689_),
    .A2(_04792_),
    .B(_04798_),
    .ZN(_01396_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09614_ (.A1(\u_cpu.rf_ram.memory[0][6] ),
    .A2(_04792_),
    .ZN(_04799_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09615_ (.A1(_02691_),
    .A2(_04792_),
    .B(_04799_),
    .ZN(_01397_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09616_ (.A1(\u_cpu.rf_ram.memory[0][7] ),
    .A2(_04792_),
    .ZN(_04800_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09617_ (.A1(_02693_),
    .A2(_04792_),
    .B(_04800_),
    .ZN(_01398_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09618_ (.A1(_02619_),
    .A2(_04349_),
    .ZN(_04801_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09619_ (.I(_04801_),
    .Z(_04802_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09620_ (.A1(\u_cpu.rf_ram.memory[98][0] ),
    .A2(_04802_),
    .ZN(_04803_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09621_ (.A1(_04622_),
    .A2(_04802_),
    .B(_04803_),
    .ZN(_01399_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09622_ (.A1(\u_cpu.rf_ram.memory[98][1] ),
    .A2(_04802_),
    .ZN(_04804_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09623_ (.A1(_04626_),
    .A2(_04802_),
    .B(_04804_),
    .ZN(_01400_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09624_ (.A1(\u_cpu.rf_ram.memory[98][2] ),
    .A2(_04802_),
    .ZN(_04805_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09625_ (.A1(_04628_),
    .A2(_04802_),
    .B(_04805_),
    .ZN(_01401_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09626_ (.A1(\u_cpu.rf_ram.memory[98][3] ),
    .A2(_04802_),
    .ZN(_04806_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09627_ (.A1(_04630_),
    .A2(_04802_),
    .B(_04806_),
    .ZN(_01402_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09628_ (.A1(\u_cpu.rf_ram.memory[98][4] ),
    .A2(_04802_),
    .ZN(_04807_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09629_ (.A1(_04632_),
    .A2(_04802_),
    .B(_04807_),
    .ZN(_01403_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09630_ (.A1(\u_cpu.rf_ram.memory[98][5] ),
    .A2(_04802_),
    .ZN(_04808_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09631_ (.A1(_04634_),
    .A2(_04802_),
    .B(_04808_),
    .ZN(_01404_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09632_ (.A1(\u_cpu.rf_ram.memory[98][6] ),
    .A2(_04802_),
    .ZN(_04809_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09633_ (.A1(_04636_),
    .A2(_04802_),
    .B(_04809_),
    .ZN(_01405_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09634_ (.A1(\u_cpu.rf_ram.memory[98][7] ),
    .A2(_04802_),
    .ZN(_04810_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09635_ (.A1(_04638_),
    .A2(_04802_),
    .B(_04810_),
    .ZN(_01406_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09636_ (.A1(_02717_),
    .A2(_04349_),
    .ZN(_04811_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09637_ (.I(_04811_),
    .Z(_04812_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09638_ (.A1(\u_cpu.rf_ram.memory[100][0] ),
    .A2(_04812_),
    .ZN(_04813_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09639_ (.A1(_04622_),
    .A2(_04812_),
    .B(_04813_),
    .ZN(_01407_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09640_ (.A1(\u_cpu.rf_ram.memory[100][1] ),
    .A2(_04812_),
    .ZN(_04814_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09641_ (.A1(_04626_),
    .A2(_04812_),
    .B(_04814_),
    .ZN(_01408_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09642_ (.A1(\u_cpu.rf_ram.memory[100][2] ),
    .A2(_04812_),
    .ZN(_04815_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09643_ (.A1(_04628_),
    .A2(_04812_),
    .B(_04815_),
    .ZN(_01409_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09644_ (.A1(\u_cpu.rf_ram.memory[100][3] ),
    .A2(_04812_),
    .ZN(_04816_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09645_ (.A1(_04630_),
    .A2(_04812_),
    .B(_04816_),
    .ZN(_01410_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09646_ (.A1(\u_cpu.rf_ram.memory[100][4] ),
    .A2(_04812_),
    .ZN(_04817_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09647_ (.A1(_04632_),
    .A2(_04812_),
    .B(_04817_),
    .ZN(_01411_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09648_ (.A1(\u_cpu.rf_ram.memory[100][5] ),
    .A2(_04812_),
    .ZN(_04818_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09649_ (.A1(_04634_),
    .A2(_04812_),
    .B(_04818_),
    .ZN(_01412_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09650_ (.A1(\u_cpu.rf_ram.memory[100][6] ),
    .A2(_04812_),
    .ZN(_04819_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09651_ (.A1(_04636_),
    .A2(_04812_),
    .B(_04819_),
    .ZN(_01413_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09652_ (.A1(\u_cpu.rf_ram.memory[100][7] ),
    .A2(_04812_),
    .ZN(_04820_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09653_ (.A1(_04638_),
    .A2(_04812_),
    .B(_04820_),
    .ZN(_01414_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09654_ (.A1(_02626_),
    .A2(_02838_),
    .ZN(_04821_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09655_ (.I(_04821_),
    .Z(_04822_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09656_ (.A1(\u_cpu.rf_ram.memory[89][0] ),
    .A2(_04822_),
    .ZN(_04823_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09657_ (.A1(_04622_),
    .A2(_04822_),
    .B(_04823_),
    .ZN(_01415_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09658_ (.A1(\u_cpu.rf_ram.memory[89][1] ),
    .A2(_04822_),
    .ZN(_04824_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09659_ (.A1(_04626_),
    .A2(_04822_),
    .B(_04824_),
    .ZN(_01416_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09660_ (.A1(\u_cpu.rf_ram.memory[89][2] ),
    .A2(_04822_),
    .ZN(_04825_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09661_ (.A1(_04628_),
    .A2(_04822_),
    .B(_04825_),
    .ZN(_01417_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09662_ (.A1(\u_cpu.rf_ram.memory[89][3] ),
    .A2(_04822_),
    .ZN(_04826_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09663_ (.A1(_04630_),
    .A2(_04822_),
    .B(_04826_),
    .ZN(_01418_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09664_ (.A1(\u_cpu.rf_ram.memory[89][4] ),
    .A2(_04822_),
    .ZN(_04827_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09665_ (.A1(_04632_),
    .A2(_04822_),
    .B(_04827_),
    .ZN(_01419_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09666_ (.A1(\u_cpu.rf_ram.memory[89][5] ),
    .A2(_04822_),
    .ZN(_04828_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09667_ (.A1(_04634_),
    .A2(_04822_),
    .B(_04828_),
    .ZN(_01420_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09668_ (.A1(\u_cpu.rf_ram.memory[89][6] ),
    .A2(_04822_),
    .ZN(_04829_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09669_ (.A1(_04636_),
    .A2(_04822_),
    .B(_04829_),
    .ZN(_01421_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09670_ (.A1(\u_cpu.rf_ram.memory[89][7] ),
    .A2(_04822_),
    .ZN(_04830_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09671_ (.A1(_04638_),
    .A2(_04822_),
    .B(_04830_),
    .ZN(_01422_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09672_ (.A1(_02677_),
    .A2(_02743_),
    .ZN(_04831_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09673_ (.I(_04831_),
    .Z(_04832_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09674_ (.A1(\u_cpu.rf_ram.memory[23][0] ),
    .A2(_04832_),
    .ZN(_04833_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09675_ (.A1(_04622_),
    .A2(_04832_),
    .B(_04833_),
    .ZN(_01423_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09676_ (.A1(\u_cpu.rf_ram.memory[23][1] ),
    .A2(_04832_),
    .ZN(_04834_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09677_ (.A1(_04626_),
    .A2(_04832_),
    .B(_04834_),
    .ZN(_01424_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09678_ (.A1(\u_cpu.rf_ram.memory[23][2] ),
    .A2(_04832_),
    .ZN(_04835_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09679_ (.A1(_04628_),
    .A2(_04832_),
    .B(_04835_),
    .ZN(_01425_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09680_ (.A1(\u_cpu.rf_ram.memory[23][3] ),
    .A2(_04832_),
    .ZN(_04836_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09681_ (.A1(_04630_),
    .A2(_04832_),
    .B(_04836_),
    .ZN(_01426_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09682_ (.A1(\u_cpu.rf_ram.memory[23][4] ),
    .A2(_04832_),
    .ZN(_04837_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09683_ (.A1(_04632_),
    .A2(_04832_),
    .B(_04837_),
    .ZN(_01427_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09684_ (.A1(\u_cpu.rf_ram.memory[23][5] ),
    .A2(_04832_),
    .ZN(_04838_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09685_ (.A1(_04634_),
    .A2(_04832_),
    .B(_04838_),
    .ZN(_01428_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09686_ (.A1(\u_cpu.rf_ram.memory[23][6] ),
    .A2(_04832_),
    .ZN(_04839_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09687_ (.A1(_04636_),
    .A2(_04832_),
    .B(_04839_),
    .ZN(_01429_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09688_ (.A1(\u_cpu.rf_ram.memory[23][7] ),
    .A2(_04832_),
    .ZN(_04840_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09689_ (.A1(_04638_),
    .A2(_04832_),
    .B(_04840_),
    .ZN(_01430_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09690_ (.A1(_03896_),
    .A2(_03611_),
    .ZN(_04841_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09691_ (.A1(\u_cpu.cpu.state.ibus_cyc ),
    .A2(_04841_),
    .ZN(_04842_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09692_ (.A1(_04309_),
    .A2(_04841_),
    .B(_04842_),
    .ZN(_01431_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _09693_ (.A1(_02273_),
    .A2(_02272_),
    .A3(\u_cpu.rf_ram.rdata[7] ),
    .Z(_04843_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09694_ (.I(_04843_),
    .Z(_01432_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _09695_ (.A1(_02273_),
    .A2(\u_cpu.rf_ram.rdata[7] ),
    .A3(\u_cpu.rf_ram_if.rtrig0 ),
    .Z(_04844_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09696_ (.I(_04844_),
    .Z(_01433_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09697_ (.A1(_02396_),
    .A2(\u_cpu.rf_ram_if.rreq_r ),
    .Z(_04845_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09698_ (.I(_04845_),
    .Z(_01434_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09699_ (.A1(\u_cpu.rf_ram_if.rcnt[0] ),
    .A2(\u_cpu.rf_ram_if.rcnt[1] ),
    .Z(_04846_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09700_ (.A1(_02912_),
    .A2(_04846_),
    .ZN(_04847_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09701_ (.A1(_02927_),
    .A2(_04847_),
    .ZN(_01435_));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09702_ (.D(_00096_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[82][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09703_ (.D(_00097_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[82][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09704_ (.D(_00098_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[82][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09705_ (.D(_00099_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[82][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09706_ (.D(_00100_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[82][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09707_ (.D(_00101_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[82][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09708_ (.D(_00102_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[82][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09709_ (.D(_00103_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[82][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09710_ (.D(_00104_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[21][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09711_ (.D(_00105_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[21][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09712_ (.D(_00106_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[21][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09713_ (.D(_00107_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[21][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09714_ (.D(_00108_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[21][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09715_ (.D(_00109_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[21][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09716_ (.D(_00110_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[21][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09717_ (.D(_00111_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[21][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09718_ (.D(_00112_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[81][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09719_ (.D(_00113_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[81][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09720_ (.D(_00114_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[81][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09721_ (.D(_00115_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[81][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09722_ (.D(_00116_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[81][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09723_ (.D(_00117_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[81][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09724_ (.D(_00118_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[81][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09725_ (.D(_00119_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[81][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09726_ (.D(_00120_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[18][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09727_ (.D(_00121_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[18][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09728_ (.D(_00122_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[18][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09729_ (.D(_00123_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[18][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09730_ (.D(_00124_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[18][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09731_ (.D(_00125_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[18][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09732_ (.D(_00126_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[18][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09733_ (.D(_00127_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[18][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09734_ (.D(_00128_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[20][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09735_ (.D(_00129_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[20][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09736_ (.D(_00130_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[20][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09737_ (.D(_00131_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[20][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09738_ (.D(_00132_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[20][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09739_ (.D(_00133_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[20][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09740_ (.D(_00134_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[20][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09741_ (.D(_00135_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[20][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09742_ (.D(_00136_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[1][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09743_ (.D(_00137_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[1][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09744_ (.D(_00138_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[1][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09745_ (.D(_00139_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[1][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09746_ (.D(_00140_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[1][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09747_ (.D(_00141_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[1][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09748_ (.D(_00142_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[1][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09749_ (.D(_00143_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[1][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09750_ (.D(_00144_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[7][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09751_ (.D(_00145_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[7][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09752_ (.D(_00146_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[7][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09753_ (.D(_00147_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[7][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09754_ (.D(_00148_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[7][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09755_ (.D(_00149_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[7][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09756_ (.D(_00150_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[7][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09757_ (.D(_00151_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[7][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09758_ (.D(_00152_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[80][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09759_ (.D(_00153_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[80][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09760_ (.D(_00154_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[80][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09761_ (.D(_00155_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[80][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09762_ (.D(_00156_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[80][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09763_ (.D(_00157_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[80][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09764_ (.D(_00158_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[80][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09765_ (.D(_00159_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[80][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09766_ (.D(_00160_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[78][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09767_ (.D(_00161_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[78][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09768_ (.D(_00162_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[78][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09769_ (.D(_00163_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[78][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09770_ (.D(_00164_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[78][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09771_ (.D(_00165_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[78][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09772_ (.D(_00166_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[78][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09773_ (.D(_00167_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[78][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09774_ (.D(_00168_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[42][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09775_ (.D(_00169_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[42][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09776_ (.D(_00170_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[42][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09777_ (.D(_00171_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[42][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09778_ (.D(_00172_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[42][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09779_ (.D(_00173_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[42][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09780_ (.D(_00174_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[42][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09781_ (.D(_00175_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[42][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09782_ (.D(_00176_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[46][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09783_ (.D(_00177_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[46][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09784_ (.D(_00178_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[46][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09785_ (.D(_00179_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[46][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09786_ (.D(_00180_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[46][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09787_ (.D(_00181_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[46][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09788_ (.D(_00182_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[46][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09789_ (.D(_00183_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[46][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09790_ (.D(_00184_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[45][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09791_ (.D(_00185_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[45][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09792_ (.D(_00186_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[45][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09793_ (.D(_00187_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[45][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09794_ (.D(_00188_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[45][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09795_ (.D(_00189_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[45][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09796_ (.D(_00190_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[45][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09797_ (.D(_00191_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[45][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09798_ (.D(_00192_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[44][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09799_ (.D(_00193_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[44][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09800_ (.D(_00194_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[44][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09801_ (.D(_00195_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[44][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09802_ (.D(_00196_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[44][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09803_ (.D(_00197_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[44][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09804_ (.D(_00198_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[44][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09805_ (.D(_00199_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[44][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09806_ (.D(_00200_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[51][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09807_ (.D(_00201_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[51][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09808_ (.D(_00202_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[51][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09809_ (.D(_00203_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[51][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09810_ (.D(_00204_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[51][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09811_ (.D(_00205_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[51][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09812_ (.D(_00206_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[51][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09813_ (.D(_00207_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[51][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09814_ (.D(_00208_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[41][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09815_ (.D(_00209_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[41][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09816_ (.D(_00210_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[41][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09817_ (.D(_00211_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[41][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09818_ (.D(_00212_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[41][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09819_ (.D(_00213_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[41][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09820_ (.D(_00214_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[41][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09821_ (.D(_00215_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[41][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09822_ (.D(_00216_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[43][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09823_ (.D(_00217_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[43][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09824_ (.D(_00218_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[43][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09825_ (.D(_00219_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[43][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09826_ (.D(_00220_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[43][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09827_ (.D(_00221_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[43][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09828_ (.D(_00222_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[43][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09829_ (.D(_00223_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[43][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09830_ (.D(_00224_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[48][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09831_ (.D(_00225_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[48][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09832_ (.D(_00226_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[48][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09833_ (.D(_00227_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[48][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09834_ (.D(_00228_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[48][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09835_ (.D(_00229_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[48][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09836_ (.D(_00230_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[48][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09837_ (.D(_00231_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[48][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09838_ (.D(_00232_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[47][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09839_ (.D(_00233_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[47][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09840_ (.D(_00234_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[47][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09841_ (.D(_00235_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[47][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09842_ (.D(_00236_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[47][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09843_ (.D(_00237_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[47][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09844_ (.D(_00238_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[47][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09845_ (.D(_00239_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[47][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09846_ (.D(_00240_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[50][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09847_ (.D(_00241_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[50][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09848_ (.D(_00242_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[50][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09849_ (.D(_00243_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[50][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09850_ (.D(_00244_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[50][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09851_ (.D(_00245_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[50][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09852_ (.D(_00246_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[50][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09853_ (.D(_00247_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[50][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09854_ (.D(_00248_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[4][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09855_ (.D(_00249_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[4][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09856_ (.D(_00250_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[4][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09857_ (.D(_00251_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[4][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09858_ (.D(_00252_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[4][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09859_ (.D(_00253_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[4][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09860_ (.D(_00254_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[4][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09861_ (.D(_00255_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[4][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09862_ (.D(_00256_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram_if.rreq_r ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09863_ (.D(_00257_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram_if.rcnt[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09864_ (.D(_00258_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram_if.rcnt[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09865_ (.D(_00259_),
    .CLK(io_in[4]),
    .Q(\u_cpu.raddr[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09866_ (.D(_00260_),
    .CLK(io_in[4]),
    .Q(\u_cpu.raddr[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09867_ (.D(_00261_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[16][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09868_ (.D(_00262_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[16][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09869_ (.D(_00263_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[16][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09870_ (.D(_00264_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[16][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09871_ (.D(_00265_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[16][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09872_ (.D(_00266_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[16][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09873_ (.D(_00267_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[16][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09874_ (.D(_00268_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[16][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09875_ (.D(_00269_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[17][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09876_ (.D(_00270_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[17][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09877_ (.D(_00271_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[17][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09878_ (.D(_00272_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[17][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09879_ (.D(_00273_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[17][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09880_ (.D(_00274_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[17][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09881_ (.D(_00275_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[17][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09882_ (.D(_00276_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[17][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09883_ (.D(_00277_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[40][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09884_ (.D(_00278_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[40][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09885_ (.D(_00279_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[40][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09886_ (.D(_00280_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[40][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09887_ (.D(_00281_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[40][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09888_ (.D(_00282_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[40][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09889_ (.D(_00283_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[40][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09890_ (.D(_00284_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[40][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09891_ (.D(_00285_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[119][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09892_ (.D(_00286_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[119][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09893_ (.D(_00287_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[119][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09894_ (.D(_00288_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[119][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09895_ (.D(_00289_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[119][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09896_ (.D(_00290_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[119][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09897_ (.D(_00291_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[119][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09898_ (.D(_00292_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[119][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09899_ (.D(_00293_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[129][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09900_ (.D(_00294_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[129][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09901_ (.D(_00295_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[129][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09902_ (.D(_00296_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[129][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09903_ (.D(_00297_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[129][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09904_ (.D(_00298_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[129][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09905_ (.D(_00299_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[129][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09906_ (.D(_00300_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[129][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09907_ (.D(_00301_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[139][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09908_ (.D(_00302_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[139][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09909_ (.D(_00303_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[139][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09910_ (.D(_00304_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[139][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09911_ (.D(_00305_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[139][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09912_ (.D(_00306_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[139][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09913_ (.D(_00307_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[139][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09914_ (.D(_00308_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[139][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09915_ (.D(_00309_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[77][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09916_ (.D(_00310_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[77][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09917_ (.D(_00311_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[77][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09918_ (.D(_00312_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[77][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09919_ (.D(_00313_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[77][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09920_ (.D(_00314_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[77][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09921_ (.D(_00315_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[77][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09922_ (.D(_00316_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[77][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09923_ (.D(_00317_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[74][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09924_ (.D(_00318_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[74][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09925_ (.D(_00319_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[74][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09926_ (.D(_00320_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[74][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09927_ (.D(_00321_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[74][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09928_ (.D(_00322_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[74][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09929_ (.D(_00323_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[74][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09930_ (.D(_00324_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[74][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09931_ (.D(_00325_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[76][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09932_ (.D(_00326_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[76][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09933_ (.D(_00327_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[76][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09934_ (.D(_00328_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[76][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09935_ (.D(_00329_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[76][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09936_ (.D(_00330_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[76][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09937_ (.D(_00331_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[76][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09938_ (.D(_00332_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[76][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09939_ (.D(_00333_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[75][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09940_ (.D(_00334_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[75][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09941_ (.D(_00335_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[75][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09942_ (.D(_00336_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[75][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09943_ (.D(_00337_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[75][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09944_ (.D(_00338_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[75][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09945_ (.D(_00339_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[75][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09946_ (.D(_00340_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[75][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09947_ (.D(_00341_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[6][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09948_ (.D(_00342_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[6][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09949_ (.D(_00343_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[6][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09950_ (.D(_00344_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[6][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09951_ (.D(_00345_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[6][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09952_ (.D(_00346_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[6][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09953_ (.D(_00347_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[6][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09954_ (.D(_00348_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[6][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09955_ (.D(_00349_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[68][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09956_ (.D(_00350_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[68][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09957_ (.D(_00351_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[68][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09958_ (.D(_00352_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[68][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09959_ (.D(_00353_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[68][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09960_ (.D(_00354_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[68][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09961_ (.D(_00355_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[68][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09962_ (.D(_00356_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[68][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09963_ (.D(_00357_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[67][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09964_ (.D(_00358_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[67][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09965_ (.D(_00359_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[67][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09966_ (.D(_00360_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[67][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09967_ (.D(_00361_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[67][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09968_ (.D(_00362_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[67][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09969_ (.D(_00363_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[67][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09970_ (.D(_00364_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[67][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09971_ (.D(_00365_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[66][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09972_ (.D(_00366_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[66][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09973_ (.D(_00367_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[66][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09974_ (.D(_00368_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[66][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09975_ (.D(_00369_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[66][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09976_ (.D(_00370_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[66][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09977_ (.D(_00371_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[66][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09978_ (.D(_00372_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[66][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09979_ (.D(_00373_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[65][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09980_ (.D(_00374_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[65][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09981_ (.D(_00375_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[65][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09982_ (.D(_00376_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[65][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09983_ (.D(_00377_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[65][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09984_ (.D(_00378_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[65][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09985_ (.D(_00379_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[65][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09986_ (.D(_00380_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[65][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09987_ (.D(_00381_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[64][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09988_ (.D(_00382_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[64][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09989_ (.D(_00383_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[64][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09990_ (.D(_00384_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[64][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09991_ (.D(_00385_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[64][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09992_ (.D(_00386_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[64][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09993_ (.D(_00387_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[64][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09994_ (.D(_00388_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[64][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09995_ (.D(_00389_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[29][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09996_ (.D(_00390_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[29][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09997_ (.D(_00391_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[29][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09998_ (.D(_00392_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[29][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09999_ (.D(_00393_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[29][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10000_ (.D(_00394_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[29][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10001_ (.D(_00395_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[29][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10002_ (.D(_00396_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[29][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10003_ (.D(_00397_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[63][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10004_ (.D(_00398_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[63][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10005_ (.D(_00399_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[63][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10006_ (.D(_00400_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[63][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10007_ (.D(_00401_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[63][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10008_ (.D(_00402_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[63][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10009_ (.D(_00403_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[63][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10010_ (.D(_00404_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[63][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10011_ (.D(_00405_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[62][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10012_ (.D(_00406_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[62][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10013_ (.D(_00407_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[62][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10014_ (.D(_00408_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[62][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10015_ (.D(_00409_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[62][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10016_ (.D(_00410_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[62][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10017_ (.D(_00411_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[62][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10018_ (.D(_00412_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[62][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10019_ (.D(_00413_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[61][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10020_ (.D(_00414_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[61][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10021_ (.D(_00415_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[61][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10022_ (.D(_00416_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[61][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10023_ (.D(_00417_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[61][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10024_ (.D(_00418_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[61][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10025_ (.D(_00419_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[61][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10026_ (.D(_00420_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[61][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10027_ (.D(_00421_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[60][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10028_ (.D(_00422_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[60][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10029_ (.D(_00423_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[60][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10030_ (.D(_00424_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[60][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10031_ (.D(_00425_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[60][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10032_ (.D(_00426_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[60][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10033_ (.D(_00427_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[60][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10034_ (.D(_00428_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[60][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10035_ (.D(_00429_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[19][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10036_ (.D(_00430_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[19][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10037_ (.D(_00431_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[19][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10038_ (.D(_00432_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[19][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10039_ (.D(_00433_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[19][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10040_ (.D(_00434_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[19][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10041_ (.D(_00435_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[19][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10042_ (.D(_00436_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[19][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10043_ (.D(_00437_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[5][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10044_ (.D(_00438_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[5][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10045_ (.D(_00439_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[5][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10046_ (.D(_00440_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[5][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10047_ (.D(_00441_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[5][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10048_ (.D(_00442_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[5][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10049_ (.D(_00443_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[5][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10050_ (.D(_00444_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[5][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10051_ (.D(_00445_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[58][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10052_ (.D(_00446_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[58][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10053_ (.D(_00447_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[58][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10054_ (.D(_00448_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[58][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10055_ (.D(_00449_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[58][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10056_ (.D(_00450_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[58][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10057_ (.D(_00451_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[58][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10058_ (.D(_00452_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[58][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10059_ (.D(_00453_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[57][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10060_ (.D(_00454_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[57][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10061_ (.D(_00455_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[57][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10062_ (.D(_00456_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[57][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10063_ (.D(_00457_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[57][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10064_ (.D(_00458_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[57][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10065_ (.D(_00459_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[57][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10066_ (.D(_00460_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[57][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10067_ (.D(_00461_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[56][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10068_ (.D(_00462_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[56][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10069_ (.D(_00463_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[56][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10070_ (.D(_00464_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[56][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10071_ (.D(_00465_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[56][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10072_ (.D(_00466_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[56][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10073_ (.D(_00467_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[56][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10074_ (.D(_00468_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[56][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10075_ (.D(_00469_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[55][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10076_ (.D(_00470_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[55][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10077_ (.D(_00471_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[55][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10078_ (.D(_00472_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[55][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10079_ (.D(_00473_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[55][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10080_ (.D(_00474_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[55][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10081_ (.D(_00475_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[55][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10082_ (.D(_00476_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[55][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10083_ (.D(_00477_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[54][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10084_ (.D(_00478_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[54][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10085_ (.D(_00479_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[54][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10086_ (.D(_00480_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[54][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10087_ (.D(_00481_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[54][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10088_ (.D(_00482_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[54][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10089_ (.D(_00483_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[54][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10090_ (.D(_00484_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[54][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10091_ (.D(_00485_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[53][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10092_ (.D(_00486_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[53][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10093_ (.D(_00487_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[53][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10094_ (.D(_00488_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[53][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10095_ (.D(_00489_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[53][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10096_ (.D(_00490_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[53][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10097_ (.D(_00491_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[53][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10098_ (.D(_00492_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[53][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10099_ (.D(_00493_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[52][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10100_ (.D(_00494_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[52][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10101_ (.D(_00495_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[52][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10102_ (.D(_00496_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[52][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10103_ (.D(_00497_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[52][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10104_ (.D(_00498_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[52][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10105_ (.D(_00499_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[52][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10106_ (.D(_00500_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[52][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10107_ (.D(_00501_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[9][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10108_ (.D(_00502_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[9][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10109_ (.D(_00503_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[9][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10110_ (.D(_00504_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[9][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10111_ (.D(_00505_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[9][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10112_ (.D(_00506_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[9][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10113_ (.D(_00507_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[9][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10114_ (.D(_00508_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[9][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10115_ (.D(_00509_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[15][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10116_ (.D(_00510_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[15][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10117_ (.D(_00511_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[15][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10118_ (.D(_00512_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[15][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10119_ (.D(_00513_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[15][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10120_ (.D(_00514_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[15][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10121_ (.D(_00515_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[15][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10122_ (.D(_00516_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[15][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10123_ (.D(_00000_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.rdata[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10124_ (.D(_00001_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.rdata[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10125_ (.D(_00002_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.rdata[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10126_ (.D(_00003_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.rdata[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10127_ (.D(_00004_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.rdata[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10128_ (.D(_00005_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.rdata[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10129_ (.D(_00006_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.rdata[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10130_ (.D(_00007_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.rdata[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10131_ (.D(_00517_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[142][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10132_ (.D(_00518_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[142][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10133_ (.D(_00519_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[142][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10134_ (.D(_00520_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[142][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10135_ (.D(_00521_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[142][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10136_ (.D(_00522_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[142][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10137_ (.D(_00523_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[142][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10138_ (.D(_00524_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[142][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10139_ (.D(_00525_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[141][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10140_ (.D(_00526_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[141][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10141_ (.D(_00527_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[141][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10142_ (.D(_00528_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[141][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10143_ (.D(_00529_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[141][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10144_ (.D(_00530_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[141][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10145_ (.D(_00531_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[141][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10146_ (.D(_00532_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[141][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10147_ (.D(_00533_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[140][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10148_ (.D(_00534_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[140][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10149_ (.D(_00535_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[140][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10150_ (.D(_00536_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[140][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10151_ (.D(_00537_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[140][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10152_ (.D(_00538_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[140][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10153_ (.D(_00539_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[140][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10154_ (.D(_00540_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[140][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10155_ (.D(_00541_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[13][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10156_ (.D(_00542_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[13][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10157_ (.D(_00543_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[13][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10158_ (.D(_00544_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[13][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10159_ (.D(_00545_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[13][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10160_ (.D(_00546_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[13][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10161_ (.D(_00547_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[13][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10162_ (.D(_00548_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[13][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10163_ (.D(_00549_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[72][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10164_ (.D(_00550_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[72][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10165_ (.D(_00551_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[72][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10166_ (.D(_00552_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[72][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10167_ (.D(_00553_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[72][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10168_ (.D(_00554_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[72][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10169_ (.D(_00555_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[72][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10170_ (.D(_00556_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[72][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10171_ (.D(_00557_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[73][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10172_ (.D(_00558_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[73][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10173_ (.D(_00559_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[73][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10174_ (.D(_00560_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[73][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10175_ (.D(_00561_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[73][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10176_ (.D(_00562_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[73][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10177_ (.D(_00563_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[73][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10178_ (.D(_00564_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[73][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10179_ (.D(_00565_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[71][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10180_ (.D(_00566_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[71][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10181_ (.D(_00567_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[71][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10182_ (.D(_00568_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[71][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10183_ (.D(_00569_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[71][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10184_ (.D(_00570_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[71][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10185_ (.D(_00571_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[71][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10186_ (.D(_00572_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[71][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10187_ (.D(_00573_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[70][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10188_ (.D(_00574_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[70][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10189_ (.D(_00575_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[70][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10190_ (.D(_00576_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[70][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10191_ (.D(_00577_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[70][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10192_ (.D(_00578_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[70][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10193_ (.D(_00579_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[70][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10194_ (.D(_00580_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[70][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10195_ (.D(_00581_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[143][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10196_ (.D(_00582_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[143][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10197_ (.D(_00583_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[143][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10198_ (.D(_00584_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[143][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10199_ (.D(_00585_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[143][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10200_ (.D(_00586_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[143][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10201_ (.D(_00587_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[143][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10202_ (.D(_00588_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[143][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10203_ (.D(_00589_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[14][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10204_ (.D(_00590_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[14][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10205_ (.D(_00591_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[14][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10206_ (.D(_00592_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[14][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10207_ (.D(_00593_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[14][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10208_ (.D(_00594_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[14][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10209_ (.D(_00595_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[14][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10210_ (.D(_00596_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[14][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10211_ (.D(_00597_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[138][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10212_ (.D(_00598_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[138][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10213_ (.D(_00599_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[138][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10214_ (.D(_00600_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[138][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10215_ (.D(_00601_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[138][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10216_ (.D(_00602_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[138][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10217_ (.D(_00603_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[138][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10218_ (.D(_00604_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[138][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10219_ (.D(_00605_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[39][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10220_ (.D(_00606_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[39][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10221_ (.D(_00607_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[39][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10222_ (.D(_00608_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[39][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10223_ (.D(_00609_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[39][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10224_ (.D(_00610_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[39][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10225_ (.D(_00611_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[39][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10226_ (.D(_00612_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[39][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10227_ (.D(_00613_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[137][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10228_ (.D(_00614_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[137][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10229_ (.D(_00615_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[137][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10230_ (.D(_00616_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[137][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10231_ (.D(_00617_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[137][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10232_ (.D(_00618_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[137][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10233_ (.D(_00619_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[137][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10234_ (.D(_00620_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[137][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10235_ (.D(_00621_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[49][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10236_ (.D(_00622_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[49][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10237_ (.D(_00623_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[49][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10238_ (.D(_00624_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[49][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10239_ (.D(_00625_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[49][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10240_ (.D(_00626_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[49][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10241_ (.D(_00627_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[49][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10242_ (.D(_00628_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[49][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10243_ (.D(_00629_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[136][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10244_ (.D(_00630_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[136][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10245_ (.D(_00631_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[136][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10246_ (.D(_00632_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[136][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10247_ (.D(_00633_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[136][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10248_ (.D(_00634_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[136][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10249_ (.D(_00635_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[136][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10250_ (.D(_00636_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[136][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10251_ (.D(_00637_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[135][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10252_ (.D(_00638_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[135][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10253_ (.D(_00639_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[135][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10254_ (.D(_00640_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[135][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10255_ (.D(_00641_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[135][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10256_ (.D(_00642_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[135][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10257_ (.D(_00643_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[135][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10258_ (.D(_00644_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[135][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10259_ (.D(_00645_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[134][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10260_ (.D(_00646_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[134][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10261_ (.D(_00647_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[134][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10262_ (.D(_00648_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[134][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10263_ (.D(_00649_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[134][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10264_ (.D(_00650_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[134][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10265_ (.D(_00651_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[134][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10266_ (.D(_00652_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[134][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10267_ (.D(_00653_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[133][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10268_ (.D(_00654_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[133][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10269_ (.D(_00655_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[133][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10270_ (.D(_00656_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[133][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10271_ (.D(_00657_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[133][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10272_ (.D(_00658_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[133][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10273_ (.D(_00659_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[133][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10274_ (.D(_00660_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[133][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10275_ (.D(_00661_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[132][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10276_ (.D(_00662_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[132][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10277_ (.D(_00663_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[132][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10278_ (.D(_00664_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[132][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10279_ (.D(_00665_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[132][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10280_ (.D(_00666_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[132][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10281_ (.D(_00667_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[132][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10282_ (.D(_00668_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[132][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10283_ (.D(_00669_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[131][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10284_ (.D(_00670_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[131][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10285_ (.D(_00671_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[131][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10286_ (.D(_00672_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[131][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10287_ (.D(_00673_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[131][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10288_ (.D(_00674_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[131][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10289_ (.D(_00675_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[131][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10290_ (.D(_00676_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[131][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10291_ (.D(_00677_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[130][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10292_ (.D(_00678_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[130][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10293_ (.D(_00679_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[130][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10294_ (.D(_00680_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[130][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10295_ (.D(_00681_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[130][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10296_ (.D(_00682_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[130][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10297_ (.D(_00683_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[130][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10298_ (.D(_00684_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[130][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10299_ (.D(_00685_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[12][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10300_ (.D(_00686_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[12][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10301_ (.D(_00687_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[12][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10302_ (.D(_00688_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[12][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10303_ (.D(_00689_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[12][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10304_ (.D(_00690_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[12][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10305_ (.D(_00691_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[12][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10306_ (.D(_00692_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[12][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10307_ (.D(_00693_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[22][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10308_ (.D(_00694_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[22][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10309_ (.D(_00695_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[22][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10310_ (.D(_00696_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[22][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10311_ (.D(_00697_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[22][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10312_ (.D(_00698_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[22][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10313_ (.D(_00699_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[22][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10314_ (.D(_00700_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[22][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10315_ (.D(_00701_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[128][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10316_ (.D(_00702_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[128][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10317_ (.D(_00703_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[128][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10318_ (.D(_00704_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[128][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10319_ (.D(_00705_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[128][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10320_ (.D(_00706_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[128][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10321_ (.D(_00707_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[128][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10322_ (.D(_00708_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[128][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10323_ (.D(_00709_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[127][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10324_ (.D(_00710_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[127][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10325_ (.D(_00711_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[127][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10326_ (.D(_00712_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[127][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10327_ (.D(_00713_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[127][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10328_ (.D(_00714_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[127][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10329_ (.D(_00715_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[127][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10330_ (.D(_00716_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[127][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10331_ (.D(_00717_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[126][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10332_ (.D(_00718_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[126][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10333_ (.D(_00719_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[126][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10334_ (.D(_00720_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[126][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10335_ (.D(_00721_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[126][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10336_ (.D(_00722_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[126][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10337_ (.D(_00723_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[126][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10338_ (.D(_00724_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[126][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10339_ (.D(_00725_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[125][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10340_ (.D(_00726_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[125][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10341_ (.D(_00727_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[125][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10342_ (.D(_00728_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[125][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10343_ (.D(_00729_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[125][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10344_ (.D(_00730_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[125][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10345_ (.D(_00731_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[125][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10346_ (.D(_00732_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[125][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10347_ (.D(_00733_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[124][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10348_ (.D(_00734_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[124][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10349_ (.D(_00735_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[124][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10350_ (.D(_00736_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[124][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10351_ (.D(_00737_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[124][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10352_ (.D(_00738_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[124][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10353_ (.D(_00739_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[124][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10354_ (.D(_00740_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[124][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10355_ (.D(_00015_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram_if.rdata1[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10356_ (.D(_00016_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram_if.rdata1[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10357_ (.D(_00017_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram_if.rdata1[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10358_ (.D(_00018_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram_if.rdata1[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10359_ (.D(_00019_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram_if.rdata1[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10360_ (.D(_00020_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram_if.rdata1[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10361_ (.D(_00008_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.alu.i_rs1 ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10362_ (.D(_00009_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram_if.rdata0[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10363_ (.D(_00010_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram_if.rdata0[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10364_ (.D(_00011_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram_if.rdata0[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10365_ (.D(_00012_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram_if.rdata0[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10366_ (.D(_00013_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram_if.rdata0[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10367_ (.D(_00014_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram_if.rdata0[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10368_ (.D(_00741_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[123][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10369_ (.D(_00742_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[123][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10370_ (.D(_00743_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[123][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10371_ (.D(_00744_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[123][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10372_ (.D(_00745_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[123][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10373_ (.D(_00746_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[123][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10374_ (.D(_00747_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[123][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10375_ (.D(_00748_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[123][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10376_ (.D(_00749_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[38][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10377_ (.D(_00750_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[38][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10378_ (.D(_00751_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[38][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10379_ (.D(_00752_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[38][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10380_ (.D(_00753_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[38][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10381_ (.D(_00754_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[38][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10382_ (.D(_00755_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[38][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10383_ (.D(_00756_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[38][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10384_ (.D(_00757_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[37][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10385_ (.D(_00758_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[37][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10386_ (.D(_00759_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[37][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10387_ (.D(_00760_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[37][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10388_ (.D(_00761_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[37][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10389_ (.D(_00762_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[37][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10390_ (.D(_00763_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[37][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10391_ (.D(_00764_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[37][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10392_ (.D(_00765_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[36][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10393_ (.D(_00766_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[36][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10394_ (.D(_00767_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[36][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10395_ (.D(_00768_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[36][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10396_ (.D(_00769_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[36][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10397_ (.D(_00770_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[36][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10398_ (.D(_00771_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[36][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10399_ (.D(_00772_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[36][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10400_ (.D(_00773_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.state.stage_two_req ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10401_ (.D(_00774_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.state.o_cnt[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10402_ (.D(_00775_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.mem_bytecnt[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10403_ (.D(_00776_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.mem_bytecnt[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10404_ (.D(_00777_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.state.o_cnt_r[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10405_ (.D(_00778_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.state.o_cnt_r[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10406_ (.D(_00779_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.state.o_cnt_r[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10407_ (.D(_00780_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.state.o_cnt_r[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10408_ (.D(_00781_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[91][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10409_ (.D(_00782_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[91][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10410_ (.D(_00783_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[91][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10411_ (.D(_00784_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[91][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10412_ (.D(_00785_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[91][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10413_ (.D(_00786_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[91][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10414_ (.D(_00787_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[91][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10415_ (.D(_00788_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[91][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10416_ (.D(_00789_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[90][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10417_ (.D(_00790_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[90][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10418_ (.D(_00791_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[90][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10419_ (.D(_00792_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[90][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10420_ (.D(_00793_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[90][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10421_ (.D(_00794_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[90][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10422_ (.D(_00795_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[90][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10423_ (.D(_00796_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[90][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10424_ (.D(_00797_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.state.genblk1.misalign_trap_sync_r ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10425_ (.D(_00798_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.mem_if.signbit ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10426_ (.D(_00799_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.ctrl.i_jump ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10427_ (.D(_00800_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.bufreg2.i_cnt_done ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10428_ (.D(_00801_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.state.init_done ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10429_ (.D(_00802_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[92][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10430_ (.D(_00803_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[92][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10431_ (.D(_00804_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[92][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10432_ (.D(_00805_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[92][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10433_ (.D(_00806_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[92][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10434_ (.D(_00807_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[92][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10435_ (.D(_00808_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[92][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10436_ (.D(_00809_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[92][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10437_ (.D(_00810_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[35][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10438_ (.D(_00811_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[35][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10439_ (.D(_00812_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[35][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10440_ (.D(_00813_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[35][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10441_ (.D(_00814_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[35][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10442_ (.D(_00815_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[35][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10443_ (.D(_00816_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[35][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10444_ (.D(_00817_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[35][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10445_ (.D(_00818_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[34][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10446_ (.D(_00819_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[34][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10447_ (.D(_00820_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[34][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10448_ (.D(_00821_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[34][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10449_ (.D(_00822_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[34][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10450_ (.D(_00823_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[34][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10451_ (.D(_00824_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[34][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10452_ (.D(_00825_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[34][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10453_ (.D(_00826_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[117][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10454_ (.D(_00827_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[117][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10455_ (.D(_00828_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[117][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10456_ (.D(_00829_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[117][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10457_ (.D(_00830_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[117][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10458_ (.D(_00831_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[117][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10459_ (.D(_00832_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[117][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10460_ (.D(_00833_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[117][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10461_ (.D(_00834_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[120][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10462_ (.D(_00835_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[120][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10463_ (.D(_00836_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[120][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10464_ (.D(_00837_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[120][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10465_ (.D(_00838_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[120][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10466_ (.D(_00839_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[120][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10467_ (.D(_00840_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[120][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10468_ (.D(_00841_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[120][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10469_ (.D(_00842_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[118][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10470_ (.D(_00843_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[118][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10471_ (.D(_00844_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[118][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10472_ (.D(_00845_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[118][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10473_ (.D(_00846_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[118][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10474_ (.D(_00847_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[118][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10475_ (.D(_00848_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[118][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10476_ (.D(_00849_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[118][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10477_ (.D(_00850_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[121][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10478_ (.D(_00851_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[121][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10479_ (.D(_00852_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[121][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10480_ (.D(_00853_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[121][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10481_ (.D(_00854_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[121][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10482_ (.D(_00855_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[121][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10483_ (.D(_00856_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[121][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10484_ (.D(_00857_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[121][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10485_ (.D(_00858_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[8][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10486_ (.D(_00859_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[8][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10487_ (.D(_00860_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[8][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10488_ (.D(_00861_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[8][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10489_ (.D(_00862_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[8][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10490_ (.D(_00863_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[8][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10491_ (.D(_00864_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[8][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10492_ (.D(_00865_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[8][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10493_ (.D(_00866_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[11][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10494_ (.D(_00867_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[11][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10495_ (.D(_00868_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[11][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10496_ (.D(_00869_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[11][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10497_ (.D(_00870_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[11][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10498_ (.D(_00871_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[11][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10499_ (.D(_00872_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[11][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10500_ (.D(_00873_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[11][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10501_ (.D(_00874_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[112][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10502_ (.D(_00875_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[112][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10503_ (.D(_00876_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[112][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10504_ (.D(_00877_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[112][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10505_ (.D(_00878_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[112][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10506_ (.D(_00879_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[112][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10507_ (.D(_00880_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[112][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10508_ (.D(_00881_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[112][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10509_ (.D(_00882_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[122][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10510_ (.D(_00883_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[122][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10511_ (.D(_00884_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[122][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10512_ (.D(_00885_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[122][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10513_ (.D(_00886_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[122][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10514_ (.D(_00887_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[122][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10515_ (.D(_00888_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[122][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10516_ (.D(_00889_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[122][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10517_ (.D(_00890_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[115][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10518_ (.D(_00891_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[115][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10519_ (.D(_00892_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[115][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10520_ (.D(_00893_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[115][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10521_ (.D(_00894_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[115][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10522_ (.D(_00895_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[115][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10523_ (.D(_00896_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[115][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10524_ (.D(_00897_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[115][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10525_ (.D(_00898_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[116][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10526_ (.D(_00899_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[116][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10527_ (.D(_00900_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[116][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10528_ (.D(_00901_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[116][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10529_ (.D(_00902_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[116][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10530_ (.D(_00903_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[116][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10531_ (.D(_00904_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[116][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10532_ (.D(_00905_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[116][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10533_ (.D(_00906_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[33][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10534_ (.D(_00907_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[33][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10535_ (.D(_00908_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[33][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10536_ (.D(_00909_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[33][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10537_ (.D(_00910_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[33][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10538_ (.D(_00911_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[33][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10539_ (.D(_00912_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[33][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10540_ (.D(_00913_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[33][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10541_ (.D(_00914_),
    .CLK(io_in[4]),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10542_ (.D(_00915_),
    .CLK(io_in[4]),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10543_ (.D(_00916_),
    .CLK(io_in[4]),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10544_ (.D(_00917_),
    .CLK(io_in[4]),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10545_ (.D(_00918_),
    .CLK(io_in[4]),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10546_ (.D(_00919_),
    .CLK(io_in[4]),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10547_ (.D(_00920_),
    .CLK(io_in[4]),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10548_ (.D(_00921_),
    .CLK(io_in[4]),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10549_ (.D(_00922_),
    .CLK(io_in[4]),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10550_ (.D(_00923_),
    .CLK(io_in[4]),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10551_ (.D(_00924_),
    .CLK(io_in[4]),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10552_ (.D(_00925_),
    .CLK(io_in[4]),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10553_ (.D(_00926_),
    .CLK(io_in[4]),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10554_ (.D(_00927_),
    .CLK(io_in[4]),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10555_ (.D(_00928_),
    .CLK(io_in[4]),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10556_ (.D(_00929_),
    .CLK(io_in[4]),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10557_ (.D(_00930_),
    .CLK(io_in[4]),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10558_ (.D(_00931_),
    .CLK(io_in[4]),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10559_ (.D(_00932_),
    .CLK(io_in[4]),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10560_ (.D(_00933_),
    .CLK(io_in[4]),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10561_ (.D(_00934_),
    .CLK(io_in[4]),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10562_ (.D(_00935_),
    .CLK(io_in[4]),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10563_ (.D(_00936_),
    .CLK(io_in[4]),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10564_ (.D(_00937_),
    .CLK(io_in[4]),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10565_ (.D(_00938_),
    .CLK(io_in[4]),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10566_ (.D(_00939_),
    .CLK(io_in[4]),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10567_ (.D(_00940_),
    .CLK(io_in[4]),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10568_ (.D(_00941_),
    .CLK(io_in[4]),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10569_ (.D(_00942_),
    .CLK(io_in[4]),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10570_ (.D(_00943_),
    .CLK(io_in[4]),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[29] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10571_ (.D(_00944_),
    .CLK(io_in[4]),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[30] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10572_ (.D(_00945_),
    .CLK(io_in[4]),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[31] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10573_ (.D(_00946_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[113][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10574_ (.D(_00947_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[113][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10575_ (.D(_00948_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[113][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10576_ (.D(_00949_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[113][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10577_ (.D(_00950_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[113][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10578_ (.D(_00951_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[113][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10579_ (.D(_00952_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[113][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10580_ (.D(_00953_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[113][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10581_ (.D(_00954_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.decode.opcode[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10582_ (.D(_00955_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.decode.opcode[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10583_ (.D(_00956_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.decode.opcode[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10584_ (.D(_00957_),
    .CLK(io_in[4]),
    .Q(\u_arbiter.i_wb_cpu_dbus_we ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10585_ (.D(_00958_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.branch_op ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10586_ (.D(_00959_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.bne_or_bge ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10587_ (.D(_00960_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.decode.co_mem_word ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10588_ (.D(_00961_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.csr_d_sel ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10589_ (.D(_00962_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.decode.co_ebreak ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10590_ (.D(_00963_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.decode.op21 ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10591_ (.D(_00964_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.decode.op22 ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10592_ (.D(_00965_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[114][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10593_ (.D(_00966_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[114][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10594_ (.D(_00967_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[114][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10595_ (.D(_00968_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[114][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10596_ (.D(_00969_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[114][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10597_ (.D(_00970_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[114][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10598_ (.D(_00971_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[114][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10599_ (.D(_00972_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[114][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10600_ (.D(_00973_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.decode.op26 ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10601_ (.D(_00974_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.immdec.imm24_20[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10602_ (.D(_00975_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.immdec.imm24_20[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10603_ (.D(_00976_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.immdec.imm24_20[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10604_ (.D(_00977_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.immdec.imm24_20[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10605_ (.D(_00978_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.immdec.imm24_20[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10606_ (.D(_00979_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.immdec.imm30_25[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10607_ (.D(_00980_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.immdec.imm30_25[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10608_ (.D(_00981_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.immdec.imm30_25[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10609_ (.D(_00982_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.immdec.imm30_25[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10610_ (.D(_00983_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.immdec.imm30_25[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10611_ (.D(_00984_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.immdec.imm30_25[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10612_ (.D(_00985_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.immdec.imm7 ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10613_ (.D(_00986_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.immdec.imm19_12_20[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10614_ (.D(_00987_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.immdec.imm19_12_20[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10615_ (.D(_00988_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.immdec.imm19_12_20[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10616_ (.D(_00989_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.immdec.imm19_12_20[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10617_ (.D(_00990_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.csr_imm ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10618_ (.D(_00991_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.immdec.imm19_12_20[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10619_ (.D(_00992_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.immdec.imm19_12_20[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10620_ (.D(_00993_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.immdec.imm19_12_20[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10621_ (.D(_00994_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.immdec.imm19_12_20[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10622_ (.D(_00995_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.immdec.imm31 ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10623_ (.D(_00996_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.genblk3.csr.timer_irq_r ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10624_ (.D(_00997_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[32][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10625_ (.D(_00998_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[32][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10626_ (.D(_00999_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[32][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10627_ (.D(_01000_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[32][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10628_ (.D(_01001_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[32][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10629_ (.D(_01002_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[32][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10630_ (.D(_01003_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[32][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10631_ (.D(_01004_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[32][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10632_ (.D(_01005_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[31][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10633_ (.D(_01006_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[31][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10634_ (.D(_01007_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[31][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10635_ (.D(_01008_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[31][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10636_ (.D(_01009_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[31][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10637_ (.D(_01010_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[31][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10638_ (.D(_01011_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[31][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10639_ (.D(_01012_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[31][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10640_ (.D(_01013_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.alu.cmp_r ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10641_ (.D(_01014_),
    .CLK(io_in[4]),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10642_ (.D(_01015_),
    .CLK(io_in[4]),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10643_ (.D(_01016_),
    .CLK(io_in[4]),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10644_ (.D(_01017_),
    .CLK(io_in[4]),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10645_ (.D(_01018_),
    .CLK(io_in[4]),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10646_ (.D(_01019_),
    .CLK(io_in[4]),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10647_ (.D(_01020_),
    .CLK(io_in[4]),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10648_ (.D(_01021_),
    .CLK(io_in[4]),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10649_ (.D(_01022_),
    .CLK(io_in[4]),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10650_ (.D(_01023_),
    .CLK(io_in[4]),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10651_ (.D(_01024_),
    .CLK(io_in[4]),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10652_ (.D(_01025_),
    .CLK(io_in[4]),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10653_ (.D(_01026_),
    .CLK(io_in[4]),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10654_ (.D(_01027_),
    .CLK(io_in[4]),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10655_ (.D(_01028_),
    .CLK(io_in[4]),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10656_ (.D(_01029_),
    .CLK(io_in[4]),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10657_ (.D(_01030_),
    .CLK(io_in[4]),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10658_ (.D(_01031_),
    .CLK(io_in[4]),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10659_ (.D(_01032_),
    .CLK(io_in[4]),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10660_ (.D(_01033_),
    .CLK(io_in[4]),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10661_ (.D(_01034_),
    .CLK(io_in[4]),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10662_ (.D(_01035_),
    .CLK(io_in[4]),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10663_ (.D(_01036_),
    .CLK(io_in[4]),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10664_ (.D(_01037_),
    .CLK(io_in[4]),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10665_ (.D(_01038_),
    .CLK(io_in[4]),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10666_ (.D(_01039_),
    .CLK(io_in[4]),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10667_ (.D(_01040_),
    .CLK(io_in[4]),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10668_ (.D(_01041_),
    .CLK(io_in[4]),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[29] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10669_ (.D(_01042_),
    .CLK(io_in[4]),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[30] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10670_ (.D(_01043_),
    .CLK(io_in[4]),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[31] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10671_ (.D(_00022_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.bufreg.c_r ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10672_ (.D(_01044_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.bufreg.lsb[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10673_ (.D(_01045_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.bufreg.lsb[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10674_ (.D(_01046_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[30][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10675_ (.D(_01047_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[30][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10676_ (.D(_01048_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[30][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10677_ (.D(_01049_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[30][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10678_ (.D(_01050_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[30][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10679_ (.D(_01051_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[30][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10680_ (.D(_01052_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[30][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10681_ (.D(_01053_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[30][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10682_ (.D(_00024_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.ctrl.pc_plus_offset_cy_r ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10683_ (.D(_00023_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.ctrl.pc_plus_4_cy_r ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10684_ (.D(_01054_),
    .CLK(io_in[4]),
    .Q(\u_arbiter.i_wb_cpu_ibus_adr[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10685_ (.D(_01055_),
    .CLK(io_in[4]),
    .Q(\u_arbiter.i_wb_cpu_ibus_adr[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10686_ (.D(_01056_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10687_ (.D(_01057_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10688_ (.D(_01058_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10689_ (.D(_01059_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10690_ (.D(_01060_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10691_ (.D(_01061_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10692_ (.D(_01062_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10693_ (.D(_01063_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10694_ (.D(_01064_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10695_ (.D(_01065_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10696_ (.D(_01066_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10697_ (.D(_01067_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10698_ (.D(_01068_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10699_ (.D(_01069_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10700_ (.D(_01070_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10701_ (.D(_01071_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10702_ (.D(_01072_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10703_ (.D(_01073_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10704_ (.D(_01074_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10705_ (.D(_01075_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10706_ (.D(_01076_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10707_ (.D(_01077_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10708_ (.D(_01078_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10709_ (.D(_01079_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10710_ (.D(_01080_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10711_ (.D(_01081_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10712_ (.D(_01082_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10713_ (.D(_01083_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[29] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10714_ (.D(_01084_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[30] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10715_ (.D(_01085_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[31] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10716_ (.D(_01086_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[109][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10717_ (.D(_01087_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[109][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10718_ (.D(_01088_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[109][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10719_ (.D(_01089_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[109][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10720_ (.D(_01090_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[109][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10721_ (.D(_01091_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[109][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10722_ (.D(_01092_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[109][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10723_ (.D(_01093_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[109][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10724_ (.D(_00021_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.alu.add_cy_r ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10725_ (.D(_01094_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[3][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10726_ (.D(_01095_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[3][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10727_ (.D(_01096_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[3][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10728_ (.D(_01097_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[3][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10729_ (.D(_01098_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[3][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10730_ (.D(_01099_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[3][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10731_ (.D(_01100_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[3][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10732_ (.D(_01101_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[3][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10733_ (.D(_01102_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[2][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10734_ (.D(_01103_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[2][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10735_ (.D(_01104_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[2][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10736_ (.D(_01105_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[2][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10737_ (.D(_01106_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[2][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10738_ (.D(_01107_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[2][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10739_ (.D(_01108_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[2][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10740_ (.D(_01109_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[2][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10741_ (.D(_01110_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[93][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10742_ (.D(_01111_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[93][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10743_ (.D(_01112_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[93][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10744_ (.D(_01113_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[93][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10745_ (.D(_01114_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[93][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10746_ (.D(_01115_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[93][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10747_ (.D(_01116_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[93][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10748_ (.D(_01117_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[93][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10749_ (.D(_01118_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.immdec.imm11_7[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10750_ (.D(_01119_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.immdec.imm11_7[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10751_ (.D(_01120_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.immdec.imm11_7[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10752_ (.D(_01121_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.immdec.imm11_7[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10753_ (.D(_01122_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.immdec.imm11_7[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10754_ (.D(_01123_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[97][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10755_ (.D(_01124_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[97][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10756_ (.D(_01125_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[97][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10757_ (.D(_01126_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[97][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10758_ (.D(_01127_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[97][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10759_ (.D(_01128_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[97][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10760_ (.D(_01129_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[97][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10761_ (.D(_01130_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[97][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10762_ (.D(_01131_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[94][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10763_ (.D(_01132_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[94][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10764_ (.D(_01133_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[94][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10765_ (.D(_01134_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[94][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10766_ (.D(_01135_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[94][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10767_ (.D(_01136_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[94][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10768_ (.D(_01137_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[94][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10769_ (.D(_01138_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[94][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10770_ (.D(_01139_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[95][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10771_ (.D(_01140_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[95][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10772_ (.D(_01141_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[95][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10773_ (.D(_01142_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[95][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10774_ (.D(_01143_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[95][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10775_ (.D(_01144_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[95][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10776_ (.D(_01145_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[95][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10777_ (.D(_01146_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[95][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10778_ (.D(_01147_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[96][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10779_ (.D(_01148_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[96][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10780_ (.D(_01149_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[96][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10781_ (.D(_01150_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[96][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10782_ (.D(_01151_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[96][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10783_ (.D(_01152_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[96][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10784_ (.D(_01153_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[96][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10785_ (.D(_01154_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[96][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10786_ (.D(_01155_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.bufreg.i_sh_signed ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10787_ (.D(_01156_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.genblk1.align.ctrl_misal ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10788_ (.D(_01157_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[28][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10789_ (.D(_01158_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[28][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10790_ (.D(_01159_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[28][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10791_ (.D(_01160_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[28][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10792_ (.D(_01161_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[28][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10793_ (.D(_01162_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[28][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10794_ (.D(_01163_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[28][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10795_ (.D(_01164_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[28][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10796_ (.D(_01165_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10797_ (.D(_01166_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10798_ (.D(_01167_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10799_ (.D(_01168_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10800_ (.D(_01169_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10801_ (.D(_01170_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10802_ (.D(_01171_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10803_ (.D(_01172_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10804_ (.D(_01173_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10805_ (.D(_01174_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10806_ (.D(_01175_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10807_ (.D(_01176_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10808_ (.D(_01177_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10809_ (.D(_01178_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10810_ (.D(_01179_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10811_ (.D(_01180_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10812_ (.D(_01181_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[101][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10813_ (.D(_01182_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[101][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10814_ (.D(_01183_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[101][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10815_ (.D(_01184_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[101][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10816_ (.D(_01185_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[101][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10817_ (.D(_01186_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[101][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10818_ (.D(_01187_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[101][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10819_ (.D(_01188_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[101][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10820_ (.D(_01189_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[102][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10821_ (.D(_01190_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[102][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10822_ (.D(_01191_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[102][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10823_ (.D(_01192_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[102][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10824_ (.D(_01193_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[102][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10825_ (.D(_01194_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[102][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10826_ (.D(_01195_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[102][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10827_ (.D(_01196_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[102][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10828_ (.D(_01197_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[103][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10829_ (.D(_01198_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[103][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10830_ (.D(_01199_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[103][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10831_ (.D(_01200_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[103][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10832_ (.D(_01201_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[103][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10833_ (.D(_01202_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[103][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10834_ (.D(_01203_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[103][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10835_ (.D(_01204_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[103][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10836_ (.D(_01205_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[104][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10837_ (.D(_01206_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[104][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10838_ (.D(_01207_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[104][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10839_ (.D(_01208_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[104][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10840_ (.D(_01209_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[104][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10841_ (.D(_01210_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[104][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10842_ (.D(_01211_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[104][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10843_ (.D(_01212_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[104][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10844_ (.D(_01213_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[99][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10845_ (.D(_01214_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[99][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10846_ (.D(_01215_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[99][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10847_ (.D(_01216_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[99][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10848_ (.D(_01217_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[99][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10849_ (.D(_01218_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[99][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10850_ (.D(_01219_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[99][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10851_ (.D(_01220_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[99][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10852_ (.D(_01221_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[79][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10853_ (.D(_01222_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[79][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10854_ (.D(_01223_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[79][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10855_ (.D(_01224_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[79][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10856_ (.D(_01225_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[79][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10857_ (.D(_01226_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[79][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10858_ (.D(_01227_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[79][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10859_ (.D(_01228_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[79][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10860_ (.D(_01229_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[105][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10861_ (.D(_01230_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[105][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10862_ (.D(_01231_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[105][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10863_ (.D(_01232_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[105][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10864_ (.D(_01233_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[105][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10865_ (.D(_01234_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[105][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10866_ (.D(_01235_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[105][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10867_ (.D(_01236_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[105][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10868_ (.D(_01237_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[106][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10869_ (.D(_01238_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[106][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10870_ (.D(_01239_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[106][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10871_ (.D(_01240_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[106][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10872_ (.D(_01241_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[106][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10873_ (.D(_01242_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[106][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10874_ (.D(_01243_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[106][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10875_ (.D(_01244_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[106][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10876_ (.D(_01245_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[107][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10877_ (.D(_01246_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[107][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10878_ (.D(_01247_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[107][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10879_ (.D(_01248_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[107][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10880_ (.D(_01249_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[107][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10881_ (.D(_01250_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[107][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10882_ (.D(_01251_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[107][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10883_ (.D(_01252_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[107][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10884_ (.D(_01253_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[83][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10885_ (.D(_01254_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[83][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10886_ (.D(_01255_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[83][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10887_ (.D(_01256_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[83][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10888_ (.D(_01257_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[83][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10889_ (.D(_01258_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[83][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10890_ (.D(_01259_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[83][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10891_ (.D(_01260_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[83][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10892_ (.D(_01261_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[108][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10893_ (.D(_01262_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[108][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10894_ (.D(_01263_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[108][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10895_ (.D(_01264_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[108][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10896_ (.D(_01265_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[108][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10897_ (.D(_01266_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[108][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10898_ (.D(_01267_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[108][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10899_ (.D(_01268_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[108][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10900_ (.D(_01269_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[69][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10901_ (.D(_01270_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[69][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10902_ (.D(_01271_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[69][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10903_ (.D(_01272_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[69][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10904_ (.D(_01273_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[69][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10905_ (.D(_01274_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[69][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10906_ (.D(_01275_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[69][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10907_ (.D(_01276_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[69][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10908_ (.D(_01277_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[84][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10909_ (.D(_01278_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[84][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10910_ (.D(_01279_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[84][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10911_ (.D(_01280_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[84][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10912_ (.D(_01281_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[84][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10913_ (.D(_01282_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[84][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10914_ (.D(_01283_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[84][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10915_ (.D(_01284_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[84][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10916_ (.D(_01285_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[59][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10917_ (.D(_01286_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[59][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10918_ (.D(_01287_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[59][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10919_ (.D(_01288_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[59][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10920_ (.D(_01289_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[59][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10921_ (.D(_01290_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[59][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10922_ (.D(_01291_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[59][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10923_ (.D(_01292_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[59][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10924_ (.D(_01293_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[10][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10925_ (.D(_01294_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[10][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10926_ (.D(_01295_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[10][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10927_ (.D(_01296_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[10][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10928_ (.D(_01297_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[10][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10929_ (.D(_01298_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[10][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10930_ (.D(_01299_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[10][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10931_ (.D(_01300_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[10][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10932_ (.D(_01301_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[85][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10933_ (.D(_01302_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[85][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10934_ (.D(_01303_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[85][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10935_ (.D(_01304_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[85][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10936_ (.D(_01305_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[85][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10937_ (.D(_01306_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[85][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10938_ (.D(_01307_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[85][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10939_ (.D(_01308_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[85][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10940_ (.D(_01309_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[110][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10941_ (.D(_01310_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[110][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10942_ (.D(_01311_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[110][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10943_ (.D(_01312_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[110][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10944_ (.D(_01313_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[110][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10945_ (.D(_01314_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[110][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10946_ (.D(_01315_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[110][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10947_ (.D(_01316_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[110][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10948_ (.D(_01317_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[86][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10949_ (.D(_01318_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[86][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10950_ (.D(_01319_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[86][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10951_ (.D(_01320_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[86][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10952_ (.D(_01321_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[86][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10953_ (.D(_01322_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[86][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10954_ (.D(_01323_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[86][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10955_ (.D(_01324_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[86][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10956_ (.D(_01325_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[111][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10957_ (.D(_01326_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[111][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10958_ (.D(_01327_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[111][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10959_ (.D(_01328_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[111][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10960_ (.D(_01329_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[111][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10961_ (.D(_01330_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[111][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10962_ (.D(_01331_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[111][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10963_ (.D(_01332_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[111][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10964_ (.D(_01333_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[87][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10965_ (.D(_01334_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[87][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10966_ (.D(_01335_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[87][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10967_ (.D(_01336_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[87][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10968_ (.D(_01337_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[87][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10969_ (.D(_01338_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[87][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10970_ (.D(_01339_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[87][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10971_ (.D(_01340_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[87][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10972_ (.D(_01341_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[88][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10973_ (.D(_01342_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[88][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10974_ (.D(_01343_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[88][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10975_ (.D(_01344_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[88][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10976_ (.D(_01345_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[88][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10977_ (.D(_01346_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[88][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10978_ (.D(_01347_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[88][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10979_ (.D(_01348_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[88][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10980_ (.D(_01349_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.genblk3.csr.mcause3_0[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10981_ (.D(_01350_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.genblk3.csr.mcause3_0[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10982_ (.D(_01351_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.genblk3.csr.mcause3_0[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10983_ (.D(_01352_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.genblk3.csr.mcause3_0[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10984_ (.D(_01353_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.genblk3.csr.mcause31 ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10985_ (.D(_01354_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.genblk3.csr.mstatus_mpie ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10986_ (.D(_01355_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.genblk3.csr.mie_mtie ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10987_ (.D(_01356_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.genblk3.csr.mstatus_mie ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10988_ (.D(_01357_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.ctrl.i_iscomp ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10989_ (.D(_01358_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.genblk3.csr.o_new_irq ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10990_ (.D(_01359_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[27][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10991_ (.D(_01360_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[27][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10992_ (.D(_01361_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[27][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10993_ (.D(_01362_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[27][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10994_ (.D(_01363_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[27][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10995_ (.D(_01364_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[27][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10996_ (.D(_01365_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[27][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10997_ (.D(_01366_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[27][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10998_ (.D(_01367_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[26][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10999_ (.D(_01368_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[26][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11000_ (.D(_01369_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[26][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11001_ (.D(_01370_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[26][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11002_ (.D(_01371_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[26][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11003_ (.D(_01372_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[26][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11004_ (.D(_01373_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[26][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11005_ (.D(_01374_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[26][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11006_ (.D(_01375_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[25][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11007_ (.D(_01376_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[25][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11008_ (.D(_01377_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[25][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11009_ (.D(_01378_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[25][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11010_ (.D(_01379_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[25][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11011_ (.D(_01380_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[25][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11012_ (.D(_01381_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[25][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11013_ (.D(_01382_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[25][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11014_ (.D(_01383_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[24][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11015_ (.D(_01384_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[24][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11016_ (.D(_01385_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[24][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11017_ (.D(_01386_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[24][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11018_ (.D(_01387_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[24][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11019_ (.D(_01388_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[24][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11020_ (.D(_01389_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[24][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11021_ (.D(_01390_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[24][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11022_ (.D(_01391_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[0][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11023_ (.D(_01392_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[0][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11024_ (.D(_01393_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[0][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11025_ (.D(_01394_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[0][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11026_ (.D(_01395_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[0][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11027_ (.D(_01396_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[0][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11028_ (.D(_01397_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[0][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11029_ (.D(_01398_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[0][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11030_ (.D(_01399_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[98][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11031_ (.D(_01400_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[98][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11032_ (.D(_01401_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[98][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11033_ (.D(_01402_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[98][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11034_ (.D(_01403_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[98][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11035_ (.D(_01404_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[98][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11036_ (.D(_01405_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[98][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11037_ (.D(_01406_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[98][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11038_ (.D(_01407_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[100][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11039_ (.D(_01408_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[100][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11040_ (.D(_01409_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[100][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11041_ (.D(_01410_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[100][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11042_ (.D(_01411_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[100][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11043_ (.D(_01412_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[100][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11044_ (.D(_01413_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[100][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11045_ (.D(_01414_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[100][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11046_ (.D(_01415_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[89][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11047_ (.D(_01416_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[89][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11048_ (.D(_01417_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[89][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11049_ (.D(_01418_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[89][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11050_ (.D(_01419_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[89][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11051_ (.D(_01420_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[89][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11052_ (.D(_01421_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[89][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11053_ (.D(_01422_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[89][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11054_ (.D(_00025_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.regzero ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11055_ (.D(_01423_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[23][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11056_ (.D(_01424_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[23][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11057_ (.D(_01425_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[23][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11058_ (.D(_01426_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[23][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11059_ (.D(_01427_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[23][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11060_ (.D(_01428_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[23][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11061_ (.D(_01429_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[23][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11062_ (.D(_01430_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[23][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11063_ (.D(_01431_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.state.ibus_cyc ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11064_ (.D(\u_cpu.rf_ram_if.wdata0_r[1] ),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram_if.wdata0_r[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11065_ (.D(\u_cpu.rf_ram_if.wdata0_r[2] ),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram_if.wdata0_r[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11066_ (.D(\u_cpu.rf_ram_if.wdata0_r[3] ),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram_if.wdata0_r[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11067_ (.D(\u_cpu.rf_ram_if.wdata0_r[4] ),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram_if.wdata0_r[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11068_ (.D(\u_cpu.rf_ram_if.wdata0_r[5] ),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram_if.wdata0_r[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11069_ (.D(\u_cpu.rf_ram_if.wdata0_r[6] ),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram_if.wdata0_r[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11070_ (.D(\u_cpu.cpu.o_wdata0 ),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram_if.wdata0_r[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11071_ (.D(\u_cpu.rf_ram_if.wtrig0 ),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram_if.genblk1.wtrig0_r ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11072_ (.D(_01432_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram_if.rdata1[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11073_ (.D(_01433_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram_if.rdata0[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11074_ (.D(_01434_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram_if.rgnt ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11075_ (.D(\u_cpu.rf_ram_if.rtrig0 ),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram_if.rtrig1 ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11076_ (.D(_01435_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram_if.rcnt[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11077_ (.D(\u_cpu.rf_ram_if.wdata1_r[1] ),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram_if.wdata1_r[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11078_ (.D(\u_cpu.rf_ram_if.wdata1_r[2] ),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram_if.wdata1_r[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11079_ (.D(\u_cpu.rf_ram_if.wdata1_r[3] ),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram_if.wdata1_r[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11080_ (.D(\u_cpu.rf_ram_if.wdata1_r[4] ),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram_if.wdata1_r[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11081_ (.D(\u_cpu.rf_ram_if.wdata1_r[5] ),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram_if.wdata1_r[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11082_ (.D(\u_cpu.rf_ram_if.wdata1_r[6] ),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram_if.wdata1_r[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11083_ (.D(\u_cpu.rf_ram_if.wdata1_r[7] ),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram_if.wdata1_r[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11084_ (.D(\u_cpu.cpu.o_wdata1 ),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram_if.wdata1_r[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11085_ (.D(\u_cpu.cpu.o_wen0 ),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram_if.wen0_r ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11086_ (.D(\u_cpu.cpu.o_wen1 ),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram_if.wen1_r ));
 gf180mcu_fd_sc_mcu7t5v0__dffnq_1 _11087_ (.D(\u_scanchain_local.module_data_in[69] ),
    .CLKN(io_in[0]),
    .Q(\u_scanchain_local.data_out ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11088_ (.D(_00026_),
    .CLK(io_in[0]),
    .Q(\u_cpu.cpu.genblk3.csr.i_mtip ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11089_ (.D(_00037_),
    .CLK(io_in[0]),
    .Q(\u_arbiter.i_wb_cpu_ack ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11090_ (.D(_00048_),
    .CLK(io_in[0]),
    .Q(\u_arbiter.i_wb_cpu_rdt[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11091_ (.D(_00059_),
    .CLK(io_in[0]),
    .Q(\u_arbiter.i_wb_cpu_rdt[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11092_ (.D(_00070_),
    .CLK(io_in[0]),
    .Q(\u_arbiter.i_wb_cpu_rdt[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11093_ (.D(_00081_),
    .CLK(io_in[0]),
    .Q(\u_arbiter.i_wb_cpu_rdt[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11094_ (.D(_00092_),
    .CLK(io_in[0]),
    .Q(\u_arbiter.i_wb_cpu_rdt[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11095_ (.D(_00093_),
    .CLK(io_in[0]),
    .Q(\u_arbiter.i_wb_cpu_rdt[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11096_ (.D(_00094_),
    .CLK(io_in[0]),
    .Q(\u_arbiter.i_wb_cpu_rdt[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11097_ (.D(_00095_),
    .CLK(io_in[0]),
    .Q(\u_arbiter.i_wb_cpu_rdt[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11098_ (.D(_00027_),
    .CLK(io_in[0]),
    .Q(\u_arbiter.i_wb_cpu_rdt[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11099_ (.D(_00028_),
    .CLK(io_in[0]),
    .Q(\u_arbiter.i_wb_cpu_rdt[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11100_ (.D(_00029_),
    .CLK(io_in[0]),
    .Q(\u_arbiter.i_wb_cpu_rdt[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11101_ (.D(_00030_),
    .CLK(io_in[0]),
    .Q(\u_arbiter.i_wb_cpu_rdt[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11102_ (.D(_00031_),
    .CLK(io_in[0]),
    .Q(\u_arbiter.i_wb_cpu_rdt[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11103_ (.D(_00032_),
    .CLK(io_in[0]),
    .Q(\u_arbiter.i_wb_cpu_rdt[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11104_ (.D(_00033_),
    .CLK(io_in[0]),
    .Q(\u_arbiter.i_wb_cpu_rdt[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11105_ (.D(_00034_),
    .CLK(io_in[0]),
    .Q(\u_arbiter.i_wb_cpu_rdt[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11106_ (.D(_00035_),
    .CLK(io_in[0]),
    .Q(\u_arbiter.i_wb_cpu_rdt[16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11107_ (.D(_00036_),
    .CLK(io_in[0]),
    .Q(\u_arbiter.i_wb_cpu_rdt[17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11108_ (.D(_00038_),
    .CLK(io_in[0]),
    .Q(\u_arbiter.i_wb_cpu_rdt[18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11109_ (.D(_00039_),
    .CLK(io_in[0]),
    .Q(\u_arbiter.i_wb_cpu_rdt[19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11110_ (.D(_00040_),
    .CLK(io_in[0]),
    .Q(\u_arbiter.i_wb_cpu_rdt[20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11111_ (.D(_00041_),
    .CLK(io_in[0]),
    .Q(\u_arbiter.i_wb_cpu_rdt[21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11112_ (.D(_00042_),
    .CLK(io_in[0]),
    .Q(\u_arbiter.i_wb_cpu_rdt[22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11113_ (.D(_00043_),
    .CLK(io_in[0]),
    .Q(\u_arbiter.i_wb_cpu_rdt[23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11114_ (.D(_00044_),
    .CLK(io_in[0]),
    .Q(\u_arbiter.i_wb_cpu_rdt[24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11115_ (.D(_00045_),
    .CLK(io_in[0]),
    .Q(\u_arbiter.i_wb_cpu_rdt[25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11116_ (.D(_00046_),
    .CLK(io_in[0]),
    .Q(\u_arbiter.i_wb_cpu_rdt[26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11117_ (.D(_00047_),
    .CLK(io_in[0]),
    .Q(\u_arbiter.i_wb_cpu_rdt[27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11118_ (.D(_00049_),
    .CLK(io_in[0]),
    .Q(\u_arbiter.i_wb_cpu_rdt[28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11119_ (.D(_00050_),
    .CLK(io_in[0]),
    .Q(\u_arbiter.i_wb_cpu_rdt[29] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11120_ (.D(_00051_),
    .CLK(io_in[0]),
    .Q(\u_arbiter.i_wb_cpu_rdt[30] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11121_ (.D(_00052_),
    .CLK(io_in[0]),
    .Q(\u_arbiter.i_wb_cpu_rdt[31] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11122_ (.D(_00053_),
    .CLK(io_in[0]),
    .Q(\u_scanchain_local.module_data_in[34] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11123_ (.D(_00054_),
    .CLK(io_in[0]),
    .Q(\u_scanchain_local.module_data_in[35] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11124_ (.D(_00055_),
    .CLK(io_in[0]),
    .Q(\u_scanchain_local.module_data_in[36] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11125_ (.D(_00056_),
    .CLK(io_in[0]),
    .Q(\u_scanchain_local.module_data_in[37] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11126_ (.D(_00057_),
    .CLK(io_in[0]),
    .Q(\u_scanchain_local.module_data_in[38] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11127_ (.D(_00058_),
    .CLK(io_in[0]),
    .Q(\u_scanchain_local.module_data_in[39] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11128_ (.D(_00060_),
    .CLK(io_in[0]),
    .Q(\u_scanchain_local.module_data_in[40] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11129_ (.D(_00061_),
    .CLK(io_in[0]),
    .Q(\u_scanchain_local.module_data_in[41] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11130_ (.D(_00062_),
    .CLK(io_in[0]),
    .Q(\u_scanchain_local.module_data_in[42] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11131_ (.D(_00063_),
    .CLK(io_in[0]),
    .Q(\u_scanchain_local.module_data_in[43] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11132_ (.D(_00064_),
    .CLK(io_in[0]),
    .Q(\u_scanchain_local.module_data_in[44] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11133_ (.D(_00065_),
    .CLK(io_in[0]),
    .Q(\u_scanchain_local.module_data_in[45] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11134_ (.D(_00066_),
    .CLK(io_in[0]),
    .Q(\u_scanchain_local.module_data_in[46] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11135_ (.D(_00067_),
    .CLK(io_in[0]),
    .Q(\u_scanchain_local.module_data_in[47] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11136_ (.D(_00068_),
    .CLK(io_in[0]),
    .Q(\u_scanchain_local.module_data_in[48] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11137_ (.D(_00069_),
    .CLK(io_in[0]),
    .Q(\u_scanchain_local.module_data_in[49] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11138_ (.D(_00071_),
    .CLK(io_in[0]),
    .Q(\u_scanchain_local.module_data_in[50] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11139_ (.D(_00072_),
    .CLK(io_in[0]),
    .Q(\u_scanchain_local.module_data_in[51] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11140_ (.D(_00073_),
    .CLK(io_in[0]),
    .Q(\u_scanchain_local.module_data_in[52] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11141_ (.D(_00074_),
    .CLK(io_in[0]),
    .Q(\u_scanchain_local.module_data_in[53] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11142_ (.D(_00075_),
    .CLK(io_in[0]),
    .Q(\u_scanchain_local.module_data_in[54] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11143_ (.D(_00076_),
    .CLK(io_in[0]),
    .Q(\u_scanchain_local.module_data_in[55] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11144_ (.D(_00077_),
    .CLK(io_in[0]),
    .Q(\u_scanchain_local.module_data_in[56] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11145_ (.D(_00078_),
    .CLK(io_in[0]),
    .Q(\u_scanchain_local.module_data_in[57] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11146_ (.D(_00079_),
    .CLK(io_in[0]),
    .Q(\u_scanchain_local.module_data_in[58] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11147_ (.D(_00080_),
    .CLK(io_in[0]),
    .Q(\u_scanchain_local.module_data_in[59] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11148_ (.D(_00082_),
    .CLK(io_in[0]),
    .Q(\u_scanchain_local.module_data_in[60] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11149_ (.D(_00083_),
    .CLK(io_in[0]),
    .Q(\u_scanchain_local.module_data_in[61] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11150_ (.D(_00084_),
    .CLK(io_in[0]),
    .Q(\u_scanchain_local.module_data_in[62] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11151_ (.D(_00085_),
    .CLK(io_in[0]),
    .Q(\u_scanchain_local.module_data_in[63] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11152_ (.D(_00086_),
    .CLK(io_in[0]),
    .Q(\u_scanchain_local.module_data_in[64] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11153_ (.D(_00087_),
    .CLK(io_in[0]),
    .Q(\u_scanchain_local.module_data_in[65] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11154_ (.D(_00088_),
    .CLK(io_in[0]),
    .Q(\u_scanchain_local.module_data_in[66] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11155_ (.D(_00089_),
    .CLK(io_in[0]),
    .Q(\u_scanchain_local.module_data_in[67] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11156_ (.D(_00090_),
    .CLK(io_in[0]),
    .Q(\u_scanchain_local.module_data_in[68] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11157_ (.D(_00091_),
    .CLK(io_in[0]),
    .Q(\u_scanchain_local.module_data_in[69] ));
 gf180mcu_fd_sc_mcu7t5v0__tiel _11158_ (.ZN(io_oeb[0]));
 gf180mcu_fd_sc_mcu7t5v0__tiel _11159_ (.ZN(io_oeb[1]));
 gf180mcu_fd_sc_mcu7t5v0__tiel _11160_ (.ZN(io_oeb[2]));
 gf180mcu_fd_sc_mcu7t5v0__tiel _11161_ (.ZN(io_oeb[3]));
 gf180mcu_fd_sc_mcu7t5v0__tiel _11162_ (.ZN(io_oeb[4]));
 gf180mcu_fd_sc_mcu7t5v0__tiel _11163_ (.ZN(io_out[2]));
 gf180mcu_fd_sc_mcu7t5v0__tiel _11164_ (.ZN(io_out[3]));
 gf180mcu_fd_sc_mcu7t5v0__tiel _11165_ (.ZN(io_out[4]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11166_ (.I(io_in[0]),
    .Z(io_out[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11167_ (.I(\u_scanchain_local.data_out ),
    .Z(io_out[1]));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_0 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_6 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_7 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_8 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_9 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_10 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_11 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_12 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_13 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_14 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_15 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_16 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_17 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_18 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_19 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_20 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_21 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_22 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_23 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_24 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_25 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_26 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_27 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_28 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_29 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_30 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_31 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_32 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_33 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_34 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_35 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_36 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_37 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_38 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_39 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_40 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_41 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_42 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_43 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_44 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_45 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_46 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_47 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_48 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_49 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_50 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_51 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_52 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_53 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_54 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_55 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_56 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_57 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_58 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_59 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_60 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_61 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_62 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_63 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_64 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_65 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_66 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_67 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_68 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_69 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_70 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_71 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_72 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_73 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_74 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_75 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_76 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_77 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_78 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_79 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_80 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_81 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_82 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_83 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_84 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_85 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_86 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_87 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_88 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_89 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_90 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_91 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_92 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_93 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_94 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_95 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_96 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_97 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_98 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_99 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_100 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_101 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_102 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_103 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_104 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_105 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_106 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_107 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_108 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_109 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_110 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_111 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_112 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_113 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_114 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_115 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_116 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_117 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_118 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_119 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_120 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_121 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_122 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_123 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_124 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_125 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_126 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_127 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_128 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_129 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_130 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_131 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_132 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_133 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_134 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_135 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_136 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_137 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_138 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_139 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_140 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_141 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_142 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_143 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_144 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_145 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_146 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_147 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_148 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_149 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_150 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_151 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_152 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_153 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_154 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_155 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_156 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_157 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_158 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_159 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_160 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_161 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_162 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_163 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_164 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_165 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_166 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_167 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_168 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_169 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_170 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_171 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_172 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_173 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_174 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_175 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_176 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_177 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_178 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_179 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_180 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_181 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_182 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_183 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_184 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_185 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_186 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_187 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_188 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_189 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_190 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_191 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_192 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_193 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_194 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_195 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_196 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_197 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_198 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_199 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_200 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_201 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_202 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_203 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_204 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_205 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_206 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_207 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_208 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_209 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_210 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_211 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_212 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_213 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_214 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_215 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_216 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_217 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_218 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_219 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_220 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_221 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_222 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_223 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_224 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_225 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_226 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_227 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_228 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_229 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_230 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_231 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_232 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_233 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_234 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_235 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_236 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_237 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_238 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_239 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_240 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_241 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_242 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_243 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_244 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_245 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_246 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_247 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_248 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_249 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_250 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_251 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_252 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_253 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_254 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_255 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_256 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_257 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_258 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_259 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_260 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_261 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_262 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_263 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_264 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_265 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_266 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_267 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_268 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_269 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_270 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_271 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_272 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_273 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_274 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_275 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_276 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_277 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_278 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_279 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_280 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_281 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_282 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_283 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_284 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_285 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_286 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_287 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_288 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2788 ();
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11157__D (.I(_00091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04900__A2 (.I(_01438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04896__A2 (.I(_01438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04891__A1 (.I(_01438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04882__A1 (.I(_01438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04880__I (.I(_01438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04876__A2 (.I(_01438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04851__I (.I(_01438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08593__A1 (.I(_01439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05707__A2 (.I(_01439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04876__A1 (.I(_01439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07862__B (.I(_01441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07855__B (.I(_01441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06599__A1 (.I(_01441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05851__A1 (.I(_01441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05831__A1 (.I(_01441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05774__A1 (.I(_01441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05770__A1 (.I(_01441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05739__A2 (.I(_01441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05712__A1 (.I(_01441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05709__I (.I(_01441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05706__A1 (.I(_01441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05683__A1 (.I(_01441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04863__A1 (.I(_01441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04856__A1 (.I(_01441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07862__C (.I(_01442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07855__A2 (.I(_01442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05784__A1 (.I(_01442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05771__B (.I(_01442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05740__A1 (.I(_01442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05734__I (.I(_01442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05708__A1 (.I(_01442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05707__A1 (.I(_01442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05692__A3 (.I(_01442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04863__A3 (.I(_01442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04856__A3 (.I(_01442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09492__A2 (.I(_01443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05775__A1 (.I(_01443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04890__A2 (.I(_01443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04872__A2 (.I(_01443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04860__A1 (.I(_01443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08567__A1 (.I(_01444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08546__A1 (.I(_01444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08497__A1 (.I(_01444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07851__A1 (.I(_01444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06589__A1 (.I(_01444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05834__A1 (.I(_01444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05784__B (.I(_01444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05743__A1 (.I(_01444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05738__I (.I(_01444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05736__B (.I(_01444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05692__A1 (.I(_01444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05689__A1 (.I(_01444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04870__A1 (.I(_01444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04859__A1 (.I(_01444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06095__A1 (.I(_01445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05790__A1 (.I(_01445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05751__A1 (.I(_01445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05744__A1 (.I(_01445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05736__A1 (.I(_01445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05733__A1 (.I(_01445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05730__I (.I(_01445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05692__A2 (.I(_01445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05684__C (.I(_01445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04870__A2 (.I(_01445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04859__A2 (.I(_01445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08850__A1 (.I(_01451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08849__B (.I(_01451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04865__B (.I(_01451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04892__A2 (.I(_01452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04882__A2 (.I(_01452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04879__A2 (.I(_01452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04866__A2 (.I(_01452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06196__A1 (.I(_01460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06128__A1 (.I(_01460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06120__A1 (.I(_01460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06116__A1 (.I(_01460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05794__A1 (.I(_01460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05791__B (.I(_01460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05726__A1 (.I(_01460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04874__C (.I(_01460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05618__A1 (.I(_01463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05530__A1 (.I(_01463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05442__A1 (.I(_01463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05354__A1 (.I(_01463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05032__I (.I(_01463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04986__I (.I(_01463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04969__I (.I(_01463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04958__I (.I(_01463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04927__I (.I(_01463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04877__I (.I(_01463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05651__A1 (.I(_01464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05609__A1 (.I(_01464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05563__A1 (.I(_01464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05475__A1 (.I(_01464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05387__A1 (.I(_01464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05357__A1 (.I(_01464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05299__A1 (.I(_01464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05269__A1 (.I(_01464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05211__A1 (.I(_01464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05181__A1 (.I(_01464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05123__A1 (.I(_01464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05093__A1 (.I(_01464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05027__A1 (.I(_01464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04980__A1 (.I(_01464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04908__I (.I(_01464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04878__I (.I(_01464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05677__A1 (.I(_01465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05671__A1 (.I(_01465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05583__A1 (.I(_01465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05499__A1 (.I(_01465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05495__A1 (.I(_01465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05411__A1 (.I(_01465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05407__A1 (.I(_01465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05323__A1 (.I(_01465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05319__A1 (.I(_01465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05235__A1 (.I(_01465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05231__A1 (.I(_01465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05147__A1 (.I(_01465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05143__A1 (.I(_01465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05059__A1 (.I(_01465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05052__A1 (.I(_01465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04905__A1 (.I(_01465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05678__C (.I(_01466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05590__C (.I(_01466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05502__C (.I(_01466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05414__C (.I(_01466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05326__C (.I(_01466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05238__C (.I(_01466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05150__C (.I(_01466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05062__C (.I(_01466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04885__A1 (.I(_01466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05827__A1 (.I(_01467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05826__A2 (.I(_01467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05825__A1 (.I(_01467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05824__A2 (.I(_01467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05823__A1 (.I(_01467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05822__A2 (.I(_01467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05821__A1 (.I(_01467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05820__A2 (.I(_01467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05819__A1 (.I(_01467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05818__A2 (.I(_01467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05817__A1 (.I(_01467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05816__A2 (.I(_01467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05815__A1 (.I(_01467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05814__A2 (.I(_01467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04906__I (.I(_01467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04881__A2 (.I(_01467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05669__B (.I(_01471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05581__B (.I(_01471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05493__B (.I(_01471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05405__B (.I(_01471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05317__B (.I(_01471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05229__B (.I(_01471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05141__B (.I(_01471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05048__B (.I(_01471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04885__A2 (.I(_01471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05680__A1 (.I(_01473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05592__A1 (.I(_01473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05504__A1 (.I(_01473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05416__A1 (.I(_01473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05328__A1 (.I(_01473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05240__A1 (.I(_01473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05152__A1 (.I(_01473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05064__A1 (.I(_01473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04904__A1 (.I(_01473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09521__A1 (.I(_01477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09520__A2 (.I(_01477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09519__A1 (.I(_01477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04891__A2 (.I(_01477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05638__B (.I(_01480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05623__B (.I(_01480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05550__B (.I(_01480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05535__B (.I(_01480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05447__B (.I(_01480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05359__B (.I(_01480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05271__B (.I(_01480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05183__B (.I(_01480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05095__B (.I(_01480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05015__I (.I(_01480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04985__B (.I(_01480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04973__I (.I(_01480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04894__I (.I(_01480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05609__B (.I(_01481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05596__B (.I(_01481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05508__B (.I(_01481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05490__B (.I(_01481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05420__B (.I(_01481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05402__B (.I(_01481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05332__B (.I(_01481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05314__B (.I(_01481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05244__B (.I(_01481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05226__B (.I(_01481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05156__B (.I(_01481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05138__B (.I(_01481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05068__B (.I(_01481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05045__B (.I(_01481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04926__B (.I(_01481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04895__I (.I(_01481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05673__B (.I(_01482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05585__B (.I(_01482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05521__B (.I(_01482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05501__B (.I(_01482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05433__B (.I(_01482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05413__B (.I(_01482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05345__B (.I(_01482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05321__B (.I(_01482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05257__B (.I(_01482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05237__B (.I(_01482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05169__B (.I(_01482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05145__B (.I(_01482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05081__B (.I(_01482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05061__B (.I(_01482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04954__B (.I(_01482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04904__A2 (.I(_01482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05628__C (.I(_01485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04996__I (.I(_01485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04899__I (.I(_01485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05601__C (.I(_01486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05570__C (.I(_01486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05513__C (.I(_01486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05482__C (.I(_01486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05425__C (.I(_01486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05394__C (.I(_01486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05337__C (.I(_01486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05306__C (.I(_01486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05249__C (.I(_01486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05218__C (.I(_01486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05161__C (.I(_01486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05130__C (.I(_01486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05073__C (.I(_01486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05035__C (.I(_01486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04936__C (.I(_01486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04904__A3 (.I(_01486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04907__A1 (.I(_01487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04902__A1 (.I(_01487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04907__A2 (.I(_01488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04902__A2 (.I(_01488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05649__A1 (.I(_01490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05561__A1 (.I(_01490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05541__A1 (.I(_01490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05473__A1 (.I(_01490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05453__A1 (.I(_01490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05385__A1 (.I(_01490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05365__A1 (.I(_01490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05297__A1 (.I(_01490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05277__A1 (.I(_01490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05209__A1 (.I(_01490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05189__A1 (.I(_01490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05121__A1 (.I(_01490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05101__A1 (.I(_01490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05025__A1 (.I(_01490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04998__A1 (.I(_01490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04904__A4 (.I(_01490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05668__A1 (.I(_01492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05630__A1 (.I(_01492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05580__A1 (.I(_01492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05542__A1 (.I(_01492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05492__A1 (.I(_01492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05454__A1 (.I(_01492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05404__A1 (.I(_01492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05366__A1 (.I(_01492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05316__A1 (.I(_01492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05278__A1 (.I(_01492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05228__A1 (.I(_01492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05190__A1 (.I(_01492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05140__A1 (.I(_01492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05102__A1 (.I(_01492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05047__A1 (.I(_01492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04999__A1 (.I(_01492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05603__A1 (.I(_01493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05587__A1 (.I(_01493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05515__A1 (.I(_01493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05506__A1 (.I(_01493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05427__A1 (.I(_01493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05418__A1 (.I(_01493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05339__A1 (.I(_01493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05330__A1 (.I(_01493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05251__A1 (.I(_01493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05242__A1 (.I(_01493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05163__A1 (.I(_01493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05154__A1 (.I(_01493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05075__A1 (.I(_01493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05066__A1 (.I(_01493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04942__A1 (.I(_01493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04918__A1 (.I(_01493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06193__B (.I(_01494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06131__A1 (.I(_01494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04982__I (.I(_01494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04970__I (.I(_01494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04944__I (.I(_01494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04922__I (.I(_01494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04910__I (.I(_01494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05613__S0 (.I(_01495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05525__S0 (.I(_01495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05437__S0 (.I(_01495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05349__S0 (.I(_01495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05261__S0 (.I(_01495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05173__S0 (.I(_01495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05085__S0 (.I(_01495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05013__I (.I(_01495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04991__I (.I(_01495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04987__I (.I(_01495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04977__I (.I(_01495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04966__I (.I(_01495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04964__S0 (.I(_01495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04959__I (.I(_01495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04937__I (.I(_01495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04911__I (.I(_01495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05640__S0 (.I(_01496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05620__S0 (.I(_01496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05552__S0 (.I(_01496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05532__S0 (.I(_01496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05464__S0 (.I(_01496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05444__S0 (.I(_01496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05376__S0 (.I(_01496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05356__S0 (.I(_01496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05288__S0 (.I(_01496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05268__S0 (.I(_01496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05200__S0 (.I(_01496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05126__S0 (.I(_01496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05112__S0 (.I(_01496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05030__S0 (.I(_01496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05010__S0 (.I(_01496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04912__I (.I(_01496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05606__S0 (.I(_01497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05593__S0 (.I(_01497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05518__S0 (.I(_01497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05505__S0 (.I(_01497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05421__S0 (.I(_01497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05417__S0 (.I(_01497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05333__S0 (.I(_01497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05329__S0 (.I(_01497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05245__S0 (.I(_01497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05241__S0 (.I(_01497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05157__S0 (.I(_01497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05153__S0 (.I(_01497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05069__S0 (.I(_01497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05065__S0 (.I(_01497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04929__S0 (.I(_01497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04917__S0 (.I(_01497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06194__A1 (.I(_01498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05020__I (.I(_01498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04992__I (.I(_01498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04983__I (.I(_01498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04971__I (.I(_01498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04946__I (.I(_01498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04914__I (.I(_01498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05613__S1 (.I(_01499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05525__S1 (.I(_01499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05437__S1 (.I(_01499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05349__S1 (.I(_01499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05261__S1 (.I(_01499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05173__S1 (.I(_01499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05085__S1 (.I(_01499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05037__I (.I(_01499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05009__I (.I(_01499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04988__I (.I(_01499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04978__I (.I(_01499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04964__S1 (.I(_01499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04960__I (.I(_01499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04939__I (.I(_01499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04924__I (.I(_01499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04915__I (.I(_01499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06133__A1 (.I(_01500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05665__S1 (.I(_01500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05635__S1 (.I(_01500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05577__S1 (.I(_01500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05547__S1 (.I(_01500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05489__S1 (.I(_01500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05459__S1 (.I(_01500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05401__S1 (.I(_01500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05371__S1 (.I(_01500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05313__S1 (.I(_01500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05283__S1 (.I(_01500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05225__S1 (.I(_01500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05137__S1 (.I(_01500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05044__S1 (.I(_01500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05040__S1 (.I(_01500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04916__I (.I(_01500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05606__S1 (.I(_01501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05593__S1 (.I(_01501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05509__S1 (.I(_01501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05505__S1 (.I(_01501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05421__S1 (.I(_01501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05417__S1 (.I(_01501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05333__S1 (.I(_01501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05329__S1 (.I(_01501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05245__S1 (.I(_01501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05241__S1 (.I(_01501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05157__S1 (.I(_01501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05153__S1 (.I(_01501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05069__S1 (.I(_01501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05065__S1 (.I(_01501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04929__S1 (.I(_01501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04917__S1 (.I(_01501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04918__A2 (.I(_01502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05614__A1 (.I(_01504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05526__A1 (.I(_01504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05438__A1 (.I(_01504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05036__I (.I(_01504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05017__I (.I(_01504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05012__I (.I(_01504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04981__I (.I(_01504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04963__I (.I(_01504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04920__I (.I(_01504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05645__A1 (.I(_01505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05616__A1 (.I(_01505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05528__A1 (.I(_01505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05440__A1 (.I(_01505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05363__A1 (.I(_01505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05352__A1 (.I(_01505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05275__A1 (.I(_01505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05264__A1 (.I(_01505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05187__A1 (.I(_01505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05176__A1 (.I(_01505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05099__A1 (.I(_01505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05088__A1 (.I(_01505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04995__A1 (.I(_01505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04968__A1 (.I(_01505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04943__I (.I(_01505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04921__I (.I(_01505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05600__A1 (.I(_01506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05596__A1 (.I(_01506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05512__A1 (.I(_01506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05508__A1 (.I(_01506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05424__A1 (.I(_01506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05420__A1 (.I(_01506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05336__A1 (.I(_01506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05332__A1 (.I(_01506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05248__A1 (.I(_01506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05244__A1 (.I(_01506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05160__A1 (.I(_01506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05156__A1 (.I(_01506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05072__A1 (.I(_01506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05068__A1 (.I(_01506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04935__A1 (.I(_01506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04926__A1 (.I(_01506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05661__S0 (.I(_01507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05656__S0 (.I(_01507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05573__S0 (.I(_01507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05568__S0 (.I(_01507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05485__S0 (.I(_01507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05480__S0 (.I(_01507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05397__S0 (.I(_01507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05392__S0 (.I(_01507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05309__S0 (.I(_01507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05304__S0 (.I(_01507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05221__S0 (.I(_01507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05216__S0 (.I(_01507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05133__S0 (.I(_01507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05128__S0 (.I(_01507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05033__S0 (.I(_01507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04923__I (.I(_01507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05604__S0 (.I(_01508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05599__S0 (.I(_01508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05516__S0 (.I(_01508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05511__S0 (.I(_01508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05423__S0 (.I(_01508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05419__S0 (.I(_01508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05335__S0 (.I(_01508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05331__S0 (.I(_01508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05247__S0 (.I(_01508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05243__S0 (.I(_01508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05159__S0 (.I(_01508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05155__S0 (.I(_01508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05071__S0 (.I(_01508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05067__S0 (.I(_01508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04931__S0 (.I(_01508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04925__S0 (.I(_01508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05604__S1 (.I(_01509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05599__S1 (.I(_01509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05511__S1 (.I(_01509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05507__S1 (.I(_01509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05423__S1 (.I(_01509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05419__S1 (.I(_01509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05335__S1 (.I(_01509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05331__S1 (.I(_01509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05247__S1 (.I(_01509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05243__S1 (.I(_01509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05159__S1 (.I(_01509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05155__S1 (.I(_01509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05071__S1 (.I(_01509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05067__S1 (.I(_01509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04931__S1 (.I(_01509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04925__S1 (.I(_01509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04926__A2 (.I(_01510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05636__A1 (.I(_01512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05632__A1 (.I(_01512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05548__A1 (.I(_01512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05544__A1 (.I(_01512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05460__A1 (.I(_01512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05456__A1 (.I(_01512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05372__A1 (.I(_01512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05314__A1 (.I(_01512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05284__A1 (.I(_01512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05226__A1 (.I(_01512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05196__A1 (.I(_01512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05138__A1 (.I(_01512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05108__A1 (.I(_01512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05045__A1 (.I(_01512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05005__A1 (.I(_01512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04928__I (.I(_01512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05598__A1 (.I(_01513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05594__A1 (.I(_01513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05521__A1 (.I(_01513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05510__A1 (.I(_01513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05433__A1 (.I(_01513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05422__A1 (.I(_01513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05345__A1 (.I(_01513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05334__A1 (.I(_01513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05257__A1 (.I(_01513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05246__A1 (.I(_01513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05169__A1 (.I(_01513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05158__A1 (.I(_01513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05081__A1 (.I(_01513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05070__A1 (.I(_01513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04954__A1 (.I(_01513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04930__A1 (.I(_01513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04930__A2 (.I(_01514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04935__A2 (.I(_01516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05634__B (.I(_01518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05614__B (.I(_01518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05526__B (.I(_01518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05438__B (.I(_01518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05350__B (.I(_01518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05262__B (.I(_01518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05174__B (.I(_01518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05086__B (.I(_01518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05022__I (.I(_01518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04994__I (.I(_01518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04965__B (.I(_01518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04934__I (.I(_01518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05600__B (.I(_01519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05574__B (.I(_01519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05512__B (.I(_01519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05486__B (.I(_01519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05424__B (.I(_01519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05398__B (.I(_01519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05336__B (.I(_01519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05310__B (.I(_01519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05248__B (.I(_01519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05222__B (.I(_01519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05160__B (.I(_01519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05134__B (.I(_01519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05072__B (.I(_01519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05041__B (.I(_01519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04949__I (.I(_01519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04935__B (.I(_01519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04999__A2 (.I(_01521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05659__S0 (.I(_01522_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05595__S0 (.I(_01522_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05571__S0 (.I(_01522_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05507__S0 (.I(_01522_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05483__S0 (.I(_01522_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05395__S0 (.I(_01522_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05307__S0 (.I(_01522_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05223__S0 (.I(_01522_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05219__S0 (.I(_01522_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05135__S0 (.I(_01522_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05131__S0 (.I(_01522_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05056__I (.I(_01522_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05049__I (.I(_01522_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05042__S0 (.I(_01522_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05038__S0 (.I(_01522_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04938__I (.I(_01522_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05674__S0 (.I(_01523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05602__S0 (.I(_01523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05586__S0 (.I(_01523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05514__S0 (.I(_01523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05430__S0 (.I(_01523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05426__S0 (.I(_01523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05342__S0 (.I(_01523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05338__S0 (.I(_01523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05254__S0 (.I(_01523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05250__S0 (.I(_01523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05166__S0 (.I(_01523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05162__S0 (.I(_01523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05078__S0 (.I(_01523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05074__S0 (.I(_01523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04951__S0 (.I(_01523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04941__S0 (.I(_01523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05631__S1 (.I(_01524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05615__S1 (.I(_01524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05543__S1 (.I(_01524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05527__S1 (.I(_01524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05455__S1 (.I(_01524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05439__S1 (.I(_01524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05367__S1 (.I(_01524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05351__S1 (.I(_01524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05263__S1 (.I(_01524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05195__S1 (.I(_01524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05175__S1 (.I(_01524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05107__S1 (.I(_01524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05087__S1 (.I(_01524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05004__S1 (.I(_01524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04967__S1 (.I(_01524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04940__I (.I(_01524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05674__S1 (.I(_01525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05602__S1 (.I(_01525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05518__S1 (.I(_01525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05514__S1 (.I(_01525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05430__S1 (.I(_01525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05426__S1 (.I(_01525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05342__S1 (.I(_01525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05338__S1 (.I(_01525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05254__S1 (.I(_01525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05250__S1 (.I(_01525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05166__S1 (.I(_01525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05162__S1 (.I(_01525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05078__S1 (.I(_01525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05074__S1 (.I(_01525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04951__S1 (.I(_01525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04941__S1 (.I(_01525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04942__A2 (.I(_01526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05607__A1 (.I(_01528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05605__A1 (.I(_01528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05519__A1 (.I(_01528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05517__A1 (.I(_01528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05431__A1 (.I(_01528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05429__A1 (.I(_01528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05343__A1 (.I(_01528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05341__A1 (.I(_01528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05255__A1 (.I(_01528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05253__A1 (.I(_01528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05167__A1 (.I(_01528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05165__A1 (.I(_01528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05079__A1 (.I(_01528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05077__A1 (.I(_01528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04952__A1 (.I(_01528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04950__A1 (.I(_01528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05665__S0 (.I(_01529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05635__S0 (.I(_01529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05577__S0 (.I(_01529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05547__S0 (.I(_01529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05489__S0 (.I(_01529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05459__S0 (.I(_01529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05401__S0 (.I(_01529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05371__S0 (.I(_01529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05313__S0 (.I(_01529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05283__S0 (.I(_01529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05225__S0 (.I(_01529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05195__S0 (.I(_01529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05137__S0 (.I(_01529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05044__S0 (.I(_01529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05040__S0 (.I(_01529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04945__I (.I(_01529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05608__S0 (.I(_01530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05597__S0 (.I(_01530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05520__S0 (.I(_01530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05509__S0 (.I(_01530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05432__S0 (.I(_01530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05428__S0 (.I(_01530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05344__S0 (.I(_01530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05340__S0 (.I(_01530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05256__S0 (.I(_01530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05252__S0 (.I(_01530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05168__S0 (.I(_01530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05164__S0 (.I(_01530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05080__S0 (.I(_01530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05076__S0 (.I(_01530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04953__S0 (.I(_01530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04948__S0 (.I(_01530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05637__S1 (.I(_01531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05617__S1 (.I(_01531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05549__S1 (.I(_01531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05529__S1 (.I(_01531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05461__S1 (.I(_01531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05441__S1 (.I(_01531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05373__S1 (.I(_01531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05353__S1 (.I(_01531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05285__S1 (.I(_01531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05265__S1 (.I(_01531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05197__S1 (.I(_01531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05177__S1 (.I(_01531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05109__S1 (.I(_01531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05089__S1 (.I(_01531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05006__S1 (.I(_01531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04947__I (.I(_01531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05608__S1 (.I(_01532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05597__S1 (.I(_01532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05520__S1 (.I(_01532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05516__S1 (.I(_01532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05432__S1 (.I(_01532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05428__S1 (.I(_01532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05344__S1 (.I(_01532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05340__S1 (.I(_01532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05256__S1 (.I(_01532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05252__S1 (.I(_01532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05168__S1 (.I(_01532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05164__S1 (.I(_01532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05080__S1 (.I(_01532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05076__S1 (.I(_01532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04953__S1 (.I(_01532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04948__S1 (.I(_01532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05677__B (.I(_01534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05605__B (.I(_01534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05589__B (.I(_01534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05517__B (.I(_01534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05497__B (.I(_01534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05429__B (.I(_01534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05409__B (.I(_01534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05341__B (.I(_01534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05325__B (.I(_01534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05253__B (.I(_01534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05233__B (.I(_01534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05165__B (.I(_01534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05149__B (.I(_01534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05077__B (.I(_01534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05055__B (.I(_01534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04950__B (.I(_01534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04957__A2 (.I(_01535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04952__A2 (.I(_01536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04975__I (.I(_01540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04956__I (.I(_01540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05667__C (.I(_01541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05610__C (.I(_01541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05579__C (.I(_01541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05522__C (.I(_01541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05491__C (.I(_01541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05434__C (.I(_01541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05403__C (.I(_01541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05346__C (.I(_01541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05315__C (.I(_01541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05258__C (.I(_01541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05227__C (.I(_01541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05170__C (.I(_01541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05139__C (.I(_01541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05082__C (.I(_01541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05046__C (.I(_01541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04957__C (.I(_01541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04999__A3 (.I(_01542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05641__A1 (.I(_01543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05621__A1 (.I(_01543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05553__A1 (.I(_01543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05533__A1 (.I(_01543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05465__A1 (.I(_01543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05445__A1 (.I(_01543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05377__A1 (.I(_01543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05348__A1 (.I(_01543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05289__A1 (.I(_01543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05260__A1 (.I(_01543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05201__A1 (.I(_01543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05172__A1 (.I(_01543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05113__A1 (.I(_01543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05084__A1 (.I(_01543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05011__A1 (.I(_01543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04962__A1 (.I(_01543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05654__S0 (.I(_01544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05611__S0 (.I(_01544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05566__S0 (.I(_01544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05523__S0 (.I(_01544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05478__S0 (.I(_01544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05435__S0 (.I(_01544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05390__S0 (.I(_01544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05347__S0 (.I(_01544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05302__S0 (.I(_01544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05259__S0 (.I(_01544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05214__S0 (.I(_01544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05171__S0 (.I(_01544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05116__S0 (.I(_01544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05083__S0 (.I(_01544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05018__S0 (.I(_01544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04961__S0 (.I(_01544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05654__S1 (.I(_01545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05611__S1 (.I(_01545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05566__S1 (.I(_01545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05523__S1 (.I(_01545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05478__S1 (.I(_01545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05435__S1 (.I(_01545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05390__S1 (.I(_01545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05347__S1 (.I(_01545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05292__S1 (.I(_01545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05259__S1 (.I(_01545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05204__S1 (.I(_01545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05171__S1 (.I(_01545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05116__S1 (.I(_01545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05083__S1 (.I(_01545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05018__S1 (.I(_01545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04961__S1 (.I(_01545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05634__A1 (.I(_01548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05623__A1 (.I(_01548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05546__A1 (.I(_01548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05535__A1 (.I(_01548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05458__A1 (.I(_01548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05447__A1 (.I(_01548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05370__A1 (.I(_01548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05350__A1 (.I(_01548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05282__A1 (.I(_01548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05262__A1 (.I(_01548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05194__A1 (.I(_01548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05174__A1 (.I(_01548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05106__A1 (.I(_01548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05086__A1 (.I(_01548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05003__A1 (.I(_01548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04965__A1 (.I(_01548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04965__A2 (.I(_01549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05631__S0 (.I(_01551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05615__S0 (.I(_01551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05543__S0 (.I(_01551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05527__S0 (.I(_01551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05455__S0 (.I(_01551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05439__S0 (.I(_01551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05367__S0 (.I(_01551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05351__S0 (.I(_01551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05279__S0 (.I(_01551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05263__S0 (.I(_01551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05191__S0 (.I(_01551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05175__S0 (.I(_01551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05107__S0 (.I(_01551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05087__S0 (.I(_01551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05004__S0 (.I(_01551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04967__S0 (.I(_01551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04976__B1 (.I(_01553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05657__A1 (.I(_01554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05647__A1 (.I(_01554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05569__A1 (.I(_01554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05559__A1 (.I(_01554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05481__A1 (.I(_01554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05471__A1 (.I(_01554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05393__A1 (.I(_01554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05383__A1 (.I(_01554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05295__A1 (.I(_01554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05266__A1 (.I(_01554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05207__A1 (.I(_01554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05178__A1 (.I(_01554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05119__A1 (.I(_01554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05090__A1 (.I(_01554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05023__A1 (.I(_01554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04974__A1 (.I(_01554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05637__S0 (.I(_01555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05617__S0 (.I(_01555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05549__S0 (.I(_01555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05529__S0 (.I(_01555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05461__S0 (.I(_01555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05441__S0 (.I(_01555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05373__S0 (.I(_01555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05353__S0 (.I(_01555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05285__S0 (.I(_01555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05265__S0 (.I(_01555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05197__S0 (.I(_01555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05177__S0 (.I(_01555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05109__S0 (.I(_01555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05089__S0 (.I(_01555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05006__S0 (.I(_01555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04972__S0 (.I(_01555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05652__S1 (.I(_01556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05642__S1 (.I(_01556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05564__S1 (.I(_01556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05554__S1 (.I(_01556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05476__S1 (.I(_01556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05466__S1 (.I(_01556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05388__S1 (.I(_01556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05378__S1 (.I(_01556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05300__S1 (.I(_01556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05290__S1 (.I(_01556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05212__S1 (.I(_01556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05202__S1 (.I(_01556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05124__S1 (.I(_01556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05114__S1 (.I(_01556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05014__S1 (.I(_01556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04972__S1 (.I(_01556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05643__B (.I(_01558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05618__B (.I(_01558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05555__B (.I(_01558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05530__B (.I(_01558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05462__B (.I(_01558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05442__B (.I(_01558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05374__B (.I(_01558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05354__B (.I(_01558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05286__B (.I(_01558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05266__B (.I(_01558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05198__B (.I(_01558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05178__B (.I(_01558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05110__B (.I(_01558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05090__B (.I(_01558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05007__B (.I(_01558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04974__B (.I(_01558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05639__C (.I(_01560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05619__C (.I(_01560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05551__C (.I(_01560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05531__C (.I(_01560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05463__C (.I(_01560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05443__C (.I(_01560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05375__C (.I(_01560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05355__C (.I(_01560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05287__C (.I(_01560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05267__C (.I(_01560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05199__C (.I(_01560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05179__C (.I(_01560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05111__C (.I(_01560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05091__C (.I(_01560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05008__C (.I(_01560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04976__C (.I(_01560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04998__A2 (.I(_01561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05663__S0 (.I(_01562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05650__S0 (.I(_01562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05575__S0 (.I(_01562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05562__S0 (.I(_01562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05487__S0 (.I(_01562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05474__S0 (.I(_01562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05399__S0 (.I(_01562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05386__S0 (.I(_01562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05311__S0 (.I(_01562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05298__S0 (.I(_01562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05210__S0 (.I(_01562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05180__S0 (.I(_01562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05122__S0 (.I(_01562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05092__S0 (.I(_01562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05026__S0 (.I(_01562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04979__S0 (.I(_01562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06263__A1 (.I(_01563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05663__S1 (.I(_01563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05650__S1 (.I(_01563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05575__S1 (.I(_01563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05562__S1 (.I(_01563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05487__S1 (.I(_01563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05474__S1 (.I(_01563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05386__S1 (.I(_01563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05298__S1 (.I(_01563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05268__S1 (.I(_01563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05210__S1 (.I(_01563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05180__S1 (.I(_01563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05122__S1 (.I(_01563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05092__S1 (.I(_01563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05026__S1 (.I(_01563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04979__S1 (.I(_01563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04980__A2 (.I(_01564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05643__A1 (.I(_01566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05638__A1 (.I(_01566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05555__A1 (.I(_01566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05550__A1 (.I(_01566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05467__A1 (.I(_01566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05462__A1 (.I(_01566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05374__A1 (.I(_01566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05359__A1 (.I(_01566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05286__A1 (.I(_01566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05271__A1 (.I(_01566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05198__A1 (.I(_01566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05183__A1 (.I(_01566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05110__A1 (.I(_01566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05095__A1 (.I(_01566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05007__A1 (.I(_01566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04985__A1 (.I(_01566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05633__S0 (.I(_01567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05622__S0 (.I(_01567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05545__S0 (.I(_01567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05534__S0 (.I(_01567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05457__S0 (.I(_01567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05446__S0 (.I(_01567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05369__S0 (.I(_01567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05358__S0 (.I(_01567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05281__S0 (.I(_01567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05270__S0 (.I(_01567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05193__S0 (.I(_01567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05182__S0 (.I(_01567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05105__S0 (.I(_01567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05094__S0 (.I(_01567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05002__S0 (.I(_01567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04984__S0 (.I(_01567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05633__S1 (.I(_01568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05622__S1 (.I(_01568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05545__S1 (.I(_01568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05534__S1 (.I(_01568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05457__S1 (.I(_01568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05446__S1 (.I(_01568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05369__S1 (.I(_01568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05358__S1 (.I(_01568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05281__S1 (.I(_01568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05270__S1 (.I(_01568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05193__S1 (.I(_01568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05182__S1 (.I(_01568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05105__S1 (.I(_01568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05094__S1 (.I(_01568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05002__S1 (.I(_01568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04984__S1 (.I(_01568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04997__A2 (.I(_01570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05625__A1 (.I(_01571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05612__A1 (.I(_01571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05537__A1 (.I(_01571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05524__A1 (.I(_01571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05449__A1 (.I(_01571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05436__A1 (.I(_01571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05368__A1 (.I(_01571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05361__A1 (.I(_01571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05280__A1 (.I(_01571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05273__A1 (.I(_01571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05192__A1 (.I(_01571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05185__A1 (.I(_01571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05104__A1 (.I(_01571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05097__A1 (.I(_01571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05001__A1 (.I(_01571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04990__A1 (.I(_01571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05644__S0 (.I(_01572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05624__S0 (.I(_01572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05556__S0 (.I(_01572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05536__S0 (.I(_01572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05468__S0 (.I(_01572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05448__S0 (.I(_01572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05380__S0 (.I(_01572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05360__S0 (.I(_01572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05292__S0 (.I(_01572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05272__S0 (.I(_01572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05204__S0 (.I(_01572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05184__S0 (.I(_01572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05103__S0 (.I(_01572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05096__S0 (.I(_01572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05000__S0 (.I(_01572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04989__S0 (.I(_01572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05644__S1 (.I(_01573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05624__S1 (.I(_01573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05556__S1 (.I(_01573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05536__S1 (.I(_01573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05468__S1 (.I(_01573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05448__S1 (.I(_01573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05380__S1 (.I(_01573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05360__S1 (.I(_01573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05279__S1 (.I(_01573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05272__S1 (.I(_01573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05191__S1 (.I(_01573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05184__S1 (.I(_01573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05103__S1 (.I(_01573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05096__S1 (.I(_01573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05000__S1 (.I(_01573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04989__S1 (.I(_01573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05646__S0 (.I(_01576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05626__S0 (.I(_01576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05558__S0 (.I(_01576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05538__S0 (.I(_01576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05470__S0 (.I(_01576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05450__S0 (.I(_01576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05382__S0 (.I(_01576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05362__S0 (.I(_01576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05294__S0 (.I(_01576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05274__S0 (.I(_01576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05206__S0 (.I(_01576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05186__S0 (.I(_01576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05118__S0 (.I(_01576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05098__S0 (.I(_01576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05021__S0 (.I(_01576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04993__S0 (.I(_01576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05646__S1 (.I(_01577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05626__S1 (.I(_01577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05558__S1 (.I(_01577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05538__S1 (.I(_01577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05470__S1 (.I(_01577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05450__S1 (.I(_01577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05382__S1 (.I(_01577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05362__S1 (.I(_01577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05294__S1 (.I(_01577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05274__S1 (.I(_01577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05206__S1 (.I(_01577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05186__S1 (.I(_01577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05118__S1 (.I(_01577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05098__S1 (.I(_01577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05028__S1 (.I(_01577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04993__S1 (.I(_01577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04995__A2 (.I(_01578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05647__B (.I(_01579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05627__B (.I(_01579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05546__B (.I(_01579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05539__B (.I(_01579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05458__B (.I(_01579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05451__B (.I(_01579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05370__B (.I(_01579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05363__B (.I(_01579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05282__B (.I(_01579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05275__B (.I(_01579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05194__B (.I(_01579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05187__B (.I(_01579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05106__B (.I(_01579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05099__B (.I(_01579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05003__B (.I(_01579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04995__B (.I(_01579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05658__C (.I(_01581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05648__C (.I(_01581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05560__C (.I(_01581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05540__C (.I(_01581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05472__C (.I(_01581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05452__C (.I(_01581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05384__C (.I(_01581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05364__C (.I(_01581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05296__C (.I(_01581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05276__C (.I(_01581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05208__C (.I(_01581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05188__C (.I(_01581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05120__C (.I(_01581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05100__C (.I(_01581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05024__C (.I(_01581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04997__C (.I(_01581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04998__A3 (.I(_01582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04999__B (.I(_01583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05008__A2 (.I(_01588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05005__A2 (.I(_01589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05025__A2 (.I(_01593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05640__S1 (.I(_01594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05620__S1 (.I(_01594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05552__S1 (.I(_01594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05532__S1 (.I(_01594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05464__S1 (.I(_01594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05444__S1 (.I(_01594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05376__S1 (.I(_01594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05356__S1 (.I(_01594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05302__S1 (.I(_01594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05288__S1 (.I(_01594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05214__S1 (.I(_01594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05200__S1 (.I(_01594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05126__S1 (.I(_01594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05112__S1 (.I(_01594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05030__S1 (.I(_01594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05010__S1 (.I(_01594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05011__A2 (.I(_01595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05653__A1 (.I(_01597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05627__A1 (.I(_01597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05565__A1 (.I(_01597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05539__A1 (.I(_01597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05477__A1 (.I(_01597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05451__A1 (.I(_01597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05389__A1 (.I(_01597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05379__A1 (.I(_01597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05301__A1 (.I(_01597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05291__A1 (.I(_01597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05213__A1 (.I(_01597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05203__A1 (.I(_01597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05125__A1 (.I(_01597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05115__A1 (.I(_01597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05029__A1 (.I(_01597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05016__A1 (.I(_01597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05652__S0 (.I(_01598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05642__S0 (.I(_01598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05564__S0 (.I(_01598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05554__S0 (.I(_01598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05476__S0 (.I(_01598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05466__S0 (.I(_01598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05388__S0 (.I(_01598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05378__S0 (.I(_01598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05300__S0 (.I(_01598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05290__S0 (.I(_01598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05212__S0 (.I(_01598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05202__S0 (.I(_01598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05124__S0 (.I(_01598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05114__S0 (.I(_01598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05028__S0 (.I(_01598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05014__S0 (.I(_01598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05666__B (.I(_01600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05653__B (.I(_01600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05578__B (.I(_01600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05565__B (.I(_01600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05477__B (.I(_01600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05467__B (.I(_01600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05389__B (.I(_01600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05379__B (.I(_01600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05301__B (.I(_01600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05291__B (.I(_01600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05213__B (.I(_01600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05203__B (.I(_01600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05125__B (.I(_01600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05115__B (.I(_01600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05029__B (.I(_01600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05016__B (.I(_01600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05664__A1 (.I(_01602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05655__A1 (.I(_01602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05567__A1 (.I(_01602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05557__A1 (.I(_01602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05479__A1 (.I(_01602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05469__A1 (.I(_01602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05391__A1 (.I(_01602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05381__A1 (.I(_01602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05303__A1 (.I(_01602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05293__A1 (.I(_01602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05215__A1 (.I(_01602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05205__A1 (.I(_01602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05127__A1 (.I(_01602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05117__A1 (.I(_01602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05031__A1 (.I(_01602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05019__A1 (.I(_01602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05661__S1 (.I(_01605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05656__S1 (.I(_01605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05573__S1 (.I(_01605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05568__S1 (.I(_01605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05485__S1 (.I(_01605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05480__S1 (.I(_01605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05397__S1 (.I(_01605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05392__S1 (.I(_01605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05309__S1 (.I(_01605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05304__S1 (.I(_01605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05221__S1 (.I(_01605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05216__S1 (.I(_01605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05133__S1 (.I(_01605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05128__S1 (.I(_01605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05033__S1 (.I(_01605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05021__S1 (.I(_01605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05023__A2 (.I(_01606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05662__B (.I(_01607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05657__B (.I(_01607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05569__B (.I(_01607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05559__B (.I(_01607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05481__B (.I(_01607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05471__B (.I(_01607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05393__B (.I(_01607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05383__B (.I(_01607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05305__B (.I(_01607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05295__B (.I(_01607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05217__B (.I(_01607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05207__B (.I(_01607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05129__B (.I(_01607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05119__B (.I(_01607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05034__B (.I(_01607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05023__B (.I(_01607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05025__A3 (.I(_01609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05048__A1 (.I(_01610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05035__A2 (.I(_01614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05031__A2 (.I(_01615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05666__A1 (.I(_01617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05662__A1 (.I(_01617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05578__A1 (.I(_01617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05574__A1 (.I(_01617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05490__A1 (.I(_01617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05486__A1 (.I(_01617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05402__A1 (.I(_01617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05398__A1 (.I(_01617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05310__A1 (.I(_01617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05305__A1 (.I(_01617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05222__A1 (.I(_01617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05217__A1 (.I(_01617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05134__A1 (.I(_01617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05129__A1 (.I(_01617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05041__A1 (.I(_01617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05034__A1 (.I(_01617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05034__A2 (.I(_01618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05660__A1 (.I(_01621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05576__A1 (.I(_01621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05572__A1 (.I(_01621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05488__A1 (.I(_01621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05484__A1 (.I(_01621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05400__A1 (.I(_01621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05396__A1 (.I(_01621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05312__A1 (.I(_01621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05308__A1 (.I(_01621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05224__A1 (.I(_01621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05220__A1 (.I(_01621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05136__A1 (.I(_01621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05132__A1 (.I(_01621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05053__I (.I(_01621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05043__A1 (.I(_01621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05039__A1 (.I(_01621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05659__S1 (.I(_01622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05595__S1 (.I(_01622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05571__S1 (.I(_01622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05483__S1 (.I(_01622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05399__S1 (.I(_01622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05395__S1 (.I(_01622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05311__S1 (.I(_01622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05307__S1 (.I(_01622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05223__S1 (.I(_01622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05219__S1 (.I(_01622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05135__S1 (.I(_01622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05131__S1 (.I(_01622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05057__I (.I(_01622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05050__I (.I(_01622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05042__S1 (.I(_01622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05038__S1 (.I(_01622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05043__A2 (.I(_01627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05046__B1 (.I(_01628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05045__A2 (.I(_01629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05047__A3 (.I(_01631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05063__A1 (.I(_01633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06609__A1 (.I(_01634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06608__A1 (.I(_01634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05672__S0 (.I(_01634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05584__S0 (.I(_01634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05496__S0 (.I(_01634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05494__S0 (.I(_01634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05408__S0 (.I(_01634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05406__S0 (.I(_01634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05320__S0 (.I(_01634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05318__S0 (.I(_01634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05232__S0 (.I(_01634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05230__S0 (.I(_01634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05144__S0 (.I(_01634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05142__S0 (.I(_01634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05054__S0 (.I(_01634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05051__S0 (.I(_01634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06612__A1 (.I(_01635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05672__S1 (.I(_01635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05584__S1 (.I(_01635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05582__S1 (.I(_01635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05496__S1 (.I(_01635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05494__S1 (.I(_01635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05408__S1 (.I(_01635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05406__S1 (.I(_01635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05320__S1 (.I(_01635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05318__S1 (.I(_01635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05232__S1 (.I(_01635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05230__S1 (.I(_01635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05144__S1 (.I(_01635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05142__S1 (.I(_01635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05054__S1 (.I(_01635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05051__S1 (.I(_01635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05052__A2 (.I(_01636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05675__A1 (.I(_01638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05673__A1 (.I(_01638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05589__A1 (.I(_01638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05585__A1 (.I(_01638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05501__A1 (.I(_01638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05497__A1 (.I(_01638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05413__A1 (.I(_01638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05409__A1 (.I(_01638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05325__A1 (.I(_01638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05321__A1 (.I(_01638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05237__A1 (.I(_01638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05233__A1 (.I(_01638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05149__A1 (.I(_01638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05145__A1 (.I(_01638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05061__A1 (.I(_01638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05055__A1 (.I(_01638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05055__A2 (.I(_01639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05676__S0 (.I(_01641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05670__S0 (.I(_01641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05588__S0 (.I(_01641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05582__S0 (.I(_01641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05500__S0 (.I(_01641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05498__S0 (.I(_01641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05412__S0 (.I(_01641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05410__S0 (.I(_01641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05324__S0 (.I(_01641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05322__S0 (.I(_01641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05236__S0 (.I(_01641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05234__S0 (.I(_01641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05148__S0 (.I(_01641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05146__S0 (.I(_01641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05060__S0 (.I(_01641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05058__S0 (.I(_01641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05676__S1 (.I(_01642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05670__S1 (.I(_01642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05588__S1 (.I(_01642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05586__S1 (.I(_01642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05500__S1 (.I(_01642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05498__S1 (.I(_01642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05412__S1 (.I(_01642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05410__S1 (.I(_01642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05324__S1 (.I(_01642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05322__S1 (.I(_01642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05236__S1 (.I(_01642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05234__S1 (.I(_01642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05148__S1 (.I(_01642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05146__S1 (.I(_01642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05060__S1 (.I(_01642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05058__S1 (.I(_01642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05059__A2 (.I(_01643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05061__A2 (.I(_01645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05063__A2 (.I(_01647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05066__A2 (.I(_01649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05068__A2 (.I(_01651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05102__A2 (.I(_01657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05075__A2 (.I(_01658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05079__A2 (.I(_01662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05102__A3 (.I(_01666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05084__A2 (.I(_01667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05086__A2 (.I(_01669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05088__A2 (.I(_01671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05091__B2 (.I(_01674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05101__A2 (.I(_01675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05100__A2 (.I(_01679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05100__B2 (.I(_01683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05101__A3 (.I(_01684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05102__B (.I(_01685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05111__A2 (.I(_01690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05108__A2 (.I(_01691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05121__A2 (.I(_01695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05113__A2 (.I(_01696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05115__A2 (.I(_01698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05117__A2 (.I(_01700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05121__A3 (.I(_01704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05141__A1 (.I(_01705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05130__A2 (.I(_01709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05127__A2 (.I(_01710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05129__A2 (.I(_01712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05132__A2 (.I(_01715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05139__B1 (.I(_01720_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05140__A3 (.I(_01723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05151__A1 (.I(_01725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05145__A2 (.I(_01728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05151__A2 (.I(_01734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05156__A2 (.I(_01738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05158__A2 (.I(_01740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05160__A2 (.I(_01742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05190__A2 (.I(_01744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05163__A2 (.I(_01745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05170__A1 (.I(_01746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05170__A2 (.I(_01748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05167__A2 (.I(_01749_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05190__A3 (.I(_01753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05174__A2 (.I(_01756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05179__A2 (.I(_01757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05179__B2 (.I(_01761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05189__A2 (.I(_01762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05188__A2 (.I(_01766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05187__A2 (.I(_01769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05189__A3 (.I(_01771_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05190__B (.I(_01772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05199__A2 (.I(_01777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05196__A2 (.I(_01778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05209__A2 (.I(_01782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05203__A2 (.I(_01785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05205__A2 (.I(_01787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05209__A3 (.I(_01791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05229__A1 (.I(_01792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05211__A2 (.I(_01793_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05218__A2 (.I(_01796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05215__A2 (.I(_01797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05217__A2 (.I(_01799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05220__A2 (.I(_01802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05222__A2 (.I(_01804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05224__A2 (.I(_01806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05227__B1 (.I(_01807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05226__A2 (.I(_01808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05228__A3 (.I(_01810_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05239__A1 (.I(_01812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05233__A2 (.I(_01815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05235__A2 (.I(_01817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05237__A2 (.I(_01819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05239__A2 (.I(_01821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05242__A2 (.I(_01823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05244__A2 (.I(_01825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05246__A2 (.I(_01827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05248__A2 (.I(_01829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05278__A2 (.I(_01831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05251__A2 (.I(_01832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05253__A2 (.I(_01834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05255__A2 (.I(_01836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05257__A2 (.I(_01838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05278__A3 (.I(_01840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05267__A1 (.I(_01842_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05262__A2 (.I(_01843_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05267__A2 (.I(_01844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05277__A2 (.I(_01849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05269__A2 (.I(_01850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05276__A2 (.I(_01853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05273__A2 (.I(_01854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05275__A2 (.I(_01856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05276__B2 (.I(_01857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05277__A3 (.I(_01858_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05278__B (.I(_01859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05287__A2 (.I(_01864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05284__A2 (.I(_01865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05297__A2 (.I(_01869_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05289__A2 (.I(_01870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05293__A2 (.I(_01874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05295__A2 (.I(_01876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05297__A3 (.I(_01878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05317__A1 (.I(_01879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05299__A2 (.I(_01880_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05306__A2 (.I(_01883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05303__A2 (.I(_01884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05305__A2 (.I(_01886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05312__A2 (.I(_01893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05314__A2 (.I(_01895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05316__A3 (.I(_01897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05327__A1 (.I(_01899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05321__A2 (.I(_01902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05327__A2 (.I(_01908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05330__A2 (.I(_01910_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05332__A2 (.I(_01912_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05336__A2 (.I(_01916_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05366__A2 (.I(_01918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05339__A2 (.I(_01919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05341__A2 (.I(_01921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05343__A2 (.I(_01923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05366__A3 (.I(_01927_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05350__A2 (.I(_01930_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05352__A2 (.I(_01932_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05365__A2 (.I(_01936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05357__A2 (.I(_01937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05364__A2 (.I(_01940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05361__A2 (.I(_01941_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05364__B2 (.I(_01944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05365__A3 (.I(_01945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05366__B (.I(_01946_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05375__A2 (.I(_01951_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05372__A2 (.I(_01952_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05385__A2 (.I(_01956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05379__A2 (.I(_01959_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05381__A2 (.I(_01961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05385__A3 (.I(_01965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05405__A1 (.I(_01966_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05387__A2 (.I(_01967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05391__A2 (.I(_01971_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05393__A2 (.I(_01973_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05404__A2 (.I(_01975_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05396__A2 (.I(_01976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05403__B1 (.I(_01981_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05402__A2 (.I(_01982_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05404__A3 (.I(_01984_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05415__A1 (.I(_01986_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05407__A2 (.I(_01987_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05409__A2 (.I(_01989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05411__A2 (.I(_01991_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05413__A2 (.I(_01993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05415__A2 (.I(_01995_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05418__A2 (.I(_01997_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05420__A2 (.I(_01999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05422__A2 (.I(_02001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05454__A2 (.I(_02005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05434__A1 (.I(_02007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05429__A2 (.I(_02008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05431__A2 (.I(_02010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05433__A2 (.I(_02012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05454__A3 (.I(_02014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05436__A2 (.I(_02015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05438__A2 (.I(_02017_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05440__A2 (.I(_02019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05453__A2 (.I(_02023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05445__A2 (.I(_02024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05449__A2 (.I(_02028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05453__A3 (.I(_02032_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05454__B (.I(_02033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05463__A2 (.I(_02038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05460__A2 (.I(_02039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05473__A2 (.I(_02043_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05465__A2 (.I(_02044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05467__A2 (.I(_02046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05469__A2 (.I(_02048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05473__A3 (.I(_02052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05493__A1 (.I(_02053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05475__A2 (.I(_02054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05482__A2 (.I(_02057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05479__A2 (.I(_02058_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05481__A2 (.I(_02060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05484__A2 (.I(_02063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05486__A2 (.I(_02065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05491__B1 (.I(_02068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05490__A2 (.I(_02069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05492__A3 (.I(_02071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05503__A1 (.I(_02073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05495__A2 (.I(_02074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05497__A2 (.I(_02076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05499__A2 (.I(_02078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05501__A2 (.I(_02080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05503__A2 (.I(_02082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05508__A2 (.I(_02086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05513__B1 (.I(_02089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05542__A2 (.I(_02092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05515__A2 (.I(_02093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05517__A2 (.I(_02095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05521__A2 (.I(_02099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05542__A3 (.I(_02101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05526__A2 (.I(_02104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05528__A2 (.I(_02106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05541__A2 (.I(_02110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05533__A2 (.I(_02111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05537__A2 (.I(_02115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05539__A2 (.I(_02117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05541__A3 (.I(_02119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05542__B (.I(_02120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05551__A2 (.I(_02125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05548__A2 (.I(_02126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05561__A2 (.I(_02130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05560__A1 (.I(_02132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05560__A2 (.I(_02134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05557__A2 (.I(_02135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05559__A2 (.I(_02137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05561__A3 (.I(_02139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05581__A1 (.I(_02140_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05563__A2 (.I(_02141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05570__A2 (.I(_02144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05567__A2 (.I(_02145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05569__A2 (.I(_02147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05572__A2 (.I(_02150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05574__A2 (.I(_02152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05576__A2 (.I(_02154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05580__A3 (.I(_02158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05591__A1 (.I(_02160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05583__A2 (.I(_02161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05585__A2 (.I(_02163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05590__B1 (.I(_02166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05589__A2 (.I(_02167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05591__A2 (.I(_02169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05596__A2 (.I(_02173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05601__B1 (.I(_02176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05630__A2 (.I(_02179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05603__A2 (.I(_02180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05609__A2 (.I(_02186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05630__A3 (.I(_02188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05614__A2 (.I(_02191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05616__A2 (.I(_02193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05629__A2 (.I(_02197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05621__A2 (.I(_02198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05625__A2 (.I(_02202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05629__A3 (.I(_02206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05630__B (.I(_02207_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05639__A2 (.I(_02212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05636__A2 (.I(_02213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05649__A2 (.I(_02217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05641__A2 (.I(_02218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05648__A2 (.I(_02221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05645__A2 (.I(_02222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05649__A3 (.I(_02226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05669__A1 (.I(_02227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05651__A2 (.I(_02228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05655__A2 (.I(_02232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05657__A2 (.I(_02234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05660__A2 (.I(_02237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05662__A2 (.I(_02239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05664__A2 (.I(_02241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05666__A2 (.I(_02243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05668__A3 (.I(_02245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05679__A1 (.I(_02247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05671__A2 (.I(_02248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05673__A2 (.I(_02250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05675__A2 (.I(_02252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09488__A1 (.I(_02259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08780__A1 (.I(_02259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08568__A1 (.I(_02259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08565__A2 (.I(_02259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08460__B (.I(_02259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08133__A1 (.I(_02259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07809__A2 (.I(_02259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06110__A1 (.I(_02259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05737__A1 (.I(_02259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05722__A1 (.I(_02259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05705__A1 (.I(_02259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05704__A1 (.I(_02259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09508__A1 (.I(_02263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09487__A1 (.I(_02263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08648__A1 (.I(_02263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07807__A2 (.I(_02263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07794__A1 (.I(_02263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06596__A1 (.I(_02263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05747__A1 (.I(_02263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05746__A1 (.I(_02263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05720__A1 (.I(_02263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05694__A1 (.I(_02263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05693__A1 (.I(_02263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08929__A1 (.I(_02264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06124__B2 (.I(_02264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05690__A2 (.I(_02264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08546__A2 (.I(_02265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08498__A1 (.I(_02265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08460__A1 (.I(_02265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08325__A1 (.I(_02265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07865__A1 (.I(_02265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06118__A1 (.I(_02265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06097__A1 (.I(_02265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05790__A2 (.I(_02265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05784__C (.I(_02265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05777__A3 (.I(_02265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05752__I (.I(_02265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05743__A2 (.I(_02265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05736__A2 (.I(_02265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05689__A2 (.I(_02265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09693__A2 (.I(_02272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05813__A1 (.I(_02272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05812__A1 (.I(_02272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05810__A1 (.I(_02272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05809__A1 (.I(_02272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05807__A1 (.I(_02272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05806__A1 (.I(_02272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05804__A1 (.I(_02272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05803__A1 (.I(_02272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05801__A1 (.I(_02272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05800__A1 (.I(_02272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05798__A1 (.I(_02272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05797__A1 (.I(_02272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05699__A1 (.I(_02272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05698__A2 (.I(_02272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09695__A1 (.I(_02273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09693__A1 (.I(_02273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05811__A1 (.I(_02273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05808__A1 (.I(_02273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05805__A1 (.I(_02273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05802__A1 (.I(_02273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05799__A1 (.I(_02273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05796__A1 (.I(_02273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05697__A2 (.I(_02273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05815__A2 (.I(_02274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05699__A2 (.I(_02274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08849__A1 (.I(_02276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05724__A2 (.I(_02276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05700__I1 (.I(_02276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08246__B2 (.I(_02277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07857__A1 (.I(_02277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05771__A2 (.I(_02277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05769__A2 (.I(_02277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05701__A2 (.I(_02277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08382__A1 (.I(_02285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07860__A1 (.I(_02285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06589__A2 (.I(_02285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05779__A1 (.I(_02285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05735__A1 (.I(_02285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05711__A1 (.I(_02285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08371__A1 (.I(_02286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07864__A1 (.I(_02286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05712__B (.I(_02286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05711__A2 (.I(_02286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05724__A1 (.I(_02289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09515__A4 (.I(_02290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08422__A1 (.I(_02290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05718__A2 (.I(_02290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09515__A3 (.I(_02291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08131__C (.I(_02291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07867__A3 (.I(_02291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07802__A1 (.I(_02291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07801__A1 (.I(_02291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07800__A1 (.I(_02291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05779__B1 (.I(_02291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05748__A2 (.I(_02291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05716__A3 (.I(_02291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09488__A3 (.I(_02292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08754__B (.I(_02292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05787__B (.I(_02292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05759__A2 (.I(_02292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05723__A2 (.I(_02292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05720__B (.I(_02292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05718__A3 (.I(_02292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09516__A1 (.I(_02293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05718__A4 (.I(_02293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09521__A2 (.I(_02301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09517__A1 (.I(_02301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05726__A2 (.I(_02301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09520__B (.I(_02303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09508__B (.I(_02303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09502__A2 (.I(_02303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09487__A2 (.I(_02303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06123__A2 (.I(_02303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06122__A1 (.I(_02303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05733__A2 (.I(_02303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05728__A2 (.I(_02303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09502__C (.I(_02305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09498__A1 (.I(_02305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08640__A1 (.I(_02305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08639__A1 (.I(_02305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08497__A2 (.I(_02305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08359__A1 (.I(_02305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07865__C (.I(_02305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07851__A2 (.I(_02305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06603__A1 (.I(_02305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06098__B (.I(_02305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06094__A1 (.I(_02305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05834__A2 (.I(_02305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05793__A1 (.I(_02305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05777__A2 (.I(_02305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05768__A1 (.I(_02305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05767__A1 (.I(_02305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08131__B (.I(_02306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05860__A2 (.I(_02306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05856__I (.I(_02306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05850__A2 (.I(_02306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05847__A1 (.I(_02306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05831__B2 (.I(_02306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05781__S0 (.I(_02306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05761__A1 (.I(_02306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05742__A1 (.I(_02306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08388__A1 (.I(_02309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07860__A2 (.I(_02309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06599__A2 (.I(_02309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05774__A2 (.I(_02309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05735__A2 (.I(_02309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08343__A1 (.I(_02313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06601__A1 (.I(_02313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06118__C (.I(_02313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06099__B (.I(_02313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05777__A1 (.I(_02313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05739__A1 (.I(_02313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08567__C (.I(_02318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05793__A2 (.I(_02318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05744__A2 (.I(_02318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08640__A2 (.I(_02320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08564__A2 (.I(_02320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08547__A1 (.I(_02320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05747__A2 (.I(_02320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06100__A1 (.I(_02322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05762__A1 (.I(_02322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05749__A1 (.I(_02322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05764__A2 (.I(_02330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05756__I (.I(_02330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08849__A2 (.I(_02334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07862__A2 (.I(_02334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06099__A1 (.I(_02334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05775__B2 (.I(_02334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05766__A2 (.I(_02334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08752__S (.I(_02335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08746__S (.I(_02335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08744__S (.I(_02335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08742__S (.I(_02335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08740__S (.I(_02335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08738__S (.I(_02335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08736__S (.I(_02335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08734__S (.I(_02335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08732__S (.I(_02335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08730__S (.I(_02335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08728__S (.I(_02335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08726__S (.I(_02335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08724__S (.I(_02335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08722__S (.I(_02335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08689__I (.I(_02335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05761__A2 (.I(_02335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05775__C (.I(_02336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05765__A1 (.I(_02336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08760__I0 (.I(_02355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08756__A1 (.I(_02355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08132__A2 (.I(_02355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08131__A2 (.I(_02355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05860__B (.I(_02355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05857__A2 (.I(_02355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05852__A1 (.I(_02355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05847__A2 (.I(_02355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05831__A2 (.I(_02355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05781__S1 (.I(_02355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05782__A2 (.I(_02356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08848__I0 (.I(_02363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05791__A1 (.I(_02363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06187__I1 (.I(_02368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05795__I (.I(_02368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05817__A2 (.I(_02369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05798__A2 (.I(_02369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05819__A2 (.I(_02371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05801__A2 (.I(_02371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05821__A2 (.I(_02373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05804__A2 (.I(_02373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06052__C (.I(_02388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06031__A1 (.I(_02388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06019__A1 (.I(_02388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05942__A1 (.I(_02388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05890__I (.I(_02388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05865__I (.I(_02388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05847__B (.I(_02388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05842__I (.I(_02388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05838__A1 (.I(_02388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05829__I (.I(_02388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06084__A1 (.I(_02389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06055__A1 (.I(_02389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06053__A1 (.I(_02389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06032__A1 (.I(_02389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06020__A1 (.I(_02389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05997__A1 (.I(_02389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05996__A1 (.I(_02389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05991__A1 (.I(_02389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05957__A1 (.I(_02389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05953__A1 (.I(_02389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05949__A1 (.I(_02389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05864__A2 (.I(_02389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05863__A2 (.I(_02389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05853__A2 (.I(_02389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05848__A2 (.I(_02389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05830__A2 (.I(_02389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08952__A2 (.I(_02392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08926__A1 (.I(_02392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08688__A1 (.I(_02392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08687__A2 (.I(_02392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08564__A1 (.I(_02392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08498__B (.I(_02392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06120__B (.I(_02392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06116__B (.I(_02392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05833__A2 (.I(_02392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09527__A1 (.I(_02395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09049__A1 (.I(_02395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08782__A1 (.I(_02395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08780__B (.I(_02395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07870__A1 (.I(_02395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07853__A1 (.I(_02395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07812__A1 (.I(_02395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07809__A1 (.I(_02395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07807__A1 (.I(_02395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07804__A1 (.I(_02395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07799__A1 (.I(_02395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07795__A1 (.I(_02395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06588__A1 (.I(_02395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05836__I (.I(_02395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09697__A1 (.I(_02396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09517__B (.I(_02396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07813__A1 (.I(_02396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07810__A1 (.I(_02396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07800__B (.I(_02396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05940__A1 (.I(_02396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05837__A1 (.I(_02396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08138__A2 (.I(_02397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06600__A2 (.I(_02397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06089__A2 (.I(_02397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06088__A1 (.I(_02397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06074__A2 (.I(_02397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06072__B (.I(_02397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06059__A2 (.I(_02397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06058__B (.I(_02397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06051__A2 (.I(_02397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06030__A2 (.I(_02397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06018__A2 (.I(_02397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05995__A2 (.I(_02397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05933__A2 (.I(_02397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05838__A2 (.I(_02397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06011__B1 (.I(_02398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06007__B1 (.I(_02398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05991__B1 (.I(_02398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05970__B1 (.I(_02398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05966__B1 (.I(_02398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05957__B1 (.I(_02398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05953__B1 (.I(_02398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05949__C1 (.I(_02398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05846__A2 (.I(_02398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05839__B (.I(_02398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09498__A2 (.I(_02400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08460__A2 (.I(_02400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08358__A1 (.I(_02400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05846__A1 (.I(_02400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06092__A1 (.I(_02402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06089__C (.I(_02402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06082__A1 (.I(_02402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06079__A1 (.I(_02402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06074__B (.I(_02402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06069__A1 (.I(_02402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06062__A1 (.I(_02402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06059__C (.I(_02402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06045__A1 (.I(_02402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06042__A1 (.I(_02402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06035__A1 (.I(_02402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06023__A1 (.I(_02402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06003__A1 (.I(_02402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06000__A1 (.I(_02402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05851__A2 (.I(_02402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05844__I (.I(_02402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06075__A1 (.I(_02403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05985__A1 (.I(_02403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05982__A1 (.I(_02403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05977__A1 (.I(_02403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05962__A1 (.I(_02403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05937__A1 (.I(_02403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05932__A1 (.I(_02403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05931__A2 (.I(_02403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05930__A1 (.I(_02403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05928__A2 (.I(_02403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05927__A1 (.I(_02403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05919__A2 (.I(_02403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05918__A2 (.I(_02403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05861__A2 (.I(_02403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05858__A2 (.I(_02403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05845__A1 (.I(_02403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08612__A2 (.I(_02411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08309__A2 (.I(_02411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08275__A2 (.I(_02411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05858__A1 (.I(_02411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05858__B1 (.I(_02413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08628__A2 (.I(_02414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08271__A2 (.I(_02414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05861__A1 (.I(_02414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08635__A2 (.I(_02416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08316__A2 (.I(_02416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08161__A1 (.I(_02416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05864__A1 (.I(_02416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06011__A1 (.I(_02418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06007__A1 (.I(_02418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05970__A1 (.I(_02418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05966__A1 (.I(_02418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05888__S (.I(_02418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05886__S (.I(_02418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05884__S (.I(_02418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05882__S (.I(_02418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05880__S (.I(_02418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05878__S (.I(_02418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05876__S (.I(_02418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05874__S (.I(_02418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05872__S (.I(_02418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05870__S (.I(_02418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05868__S (.I(_02418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05866__S (.I(_02418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05924__S (.I(_02431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05922__S (.I(_02431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05920__S (.I(_02431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05915__S (.I(_02431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05913__S (.I(_02431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05911__S (.I(_02431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05909__S (.I(_02431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05907__S (.I(_02431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05905__S (.I(_02431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05903__S (.I(_02431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05901__S (.I(_02431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05899__S (.I(_02431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05897__S (.I(_02431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05895__S (.I(_02431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05893__S (.I(_02431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05891__S (.I(_02431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06078__A1 (.I(_02456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06068__B (.I(_02456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06041__A1 (.I(_02456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06012__A1 (.I(_02456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06008__A1 (.I(_02456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05990__B (.I(_02456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05981__B (.I(_02456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05976__A1 (.I(_02456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05971__A1 (.I(_02456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05967__A1 (.I(_02456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05958__A1 (.I(_02456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05954__A1 (.I(_02456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05938__A2 (.I(_02456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05935__A2 (.I(_02456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09047__A3 (.I(_02461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08267__A2 (.I(_02461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06585__A2 (.I(_02461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06050__A1 (.I(_02461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06029__A1 (.I(_02461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06017__C (.I(_02461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05993__B (.I(_02461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05961__A2 (.I(_02461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05942__A2 (.I(_02461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06093__A1 (.I(_02463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06083__A1 (.I(_02463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06063__A1 (.I(_02463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06046__A1 (.I(_02463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06036__A1 (.I(_02463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06024__A1 (.I(_02463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06004__A1 (.I(_02463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06001__A1 (.I(_02463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05986__A1 (.I(_02463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05963__A1 (.I(_02463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05949__B1 (.I(_02463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08299__A1 (.I(_02464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08297__S (.I(_02464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08296__S (.I(_02464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08295__S (.I(_02464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08294__A1 (.I(_02464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08293__A1 (.I(_02464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06584__I (.I(_02464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05959__A1 (.I(_02464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05945__I (.I(_02464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08348__A1 (.I(_02465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08319__S (.I(_02465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08316__A1 (.I(_02465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08315__A1 (.I(_02465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08313__S (.I(_02465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08312__S (.I(_02465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08288__A1 (.I(_02465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08285__A1 (.I(_02465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08279__A1 (.I(_02465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08277__S (.I(_02465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08275__A1 (.I(_02465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08274__A1 (.I(_02465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08272__S (.I(_02465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08271__A1 (.I(_02465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08270__A1 (.I(_02465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05946__I (.I(_02465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08594__S (.I(_02466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08512__S (.I(_02466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08470__S (.I(_02466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08441__S (.I(_02466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08412__S (.I(_02466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08378__S (.I(_02466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08373__A1 (.I(_02466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08354__A1 (.I(_02466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08347__S (.I(_02466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08331__A1 (.I(_02466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08317__S (.I(_02466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08310__A1 (.I(_02466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08309__A1 (.I(_02466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08306__A1 (.I(_02466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08304__S (.I(_02466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05947__I (.I(_02466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09048__A1 (.I(_02467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08643__S (.I(_02467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08636__A1 (.I(_02467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08635__A1 (.I(_02467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08628__A1 (.I(_02467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08627__A1 (.I(_02467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08538__S (.I(_02467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08532__S (.I(_02467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08525__S (.I(_02467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08496__S (.I(_02467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08484__S (.I(_02467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08401__S (.I(_02467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08390__S (.I(_02467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05955__A1 (.I(_02467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05951__A1 (.I(_02467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05948__A1 (.I(_02467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06092__B1 (.I(_02478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06082__B1 (.I(_02478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06079__B1 (.I(_02478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06069__B1 (.I(_02478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06062__B1 (.I(_02478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06045__B1 (.I(_02478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06042__B1 (.I(_02478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06035__B1 (.I(_02478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06023__B1 (.I(_02478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06003__B1 (.I(_02478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06000__B1 (.I(_02478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05985__B1 (.I(_02478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05982__B1 (.I(_02478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05977__B1 (.I(_02478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05962__B1 (.I(_02478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05988__A3 (.I(_02487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05980__A3 (.I(_02487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05975__A2 (.I(_02487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05974__A2 (.I(_02487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06016__A3 (.I(_02499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05999__A3 (.I(_02499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05998__A2 (.I(_02499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05994__A2 (.I(_02499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05993__A2 (.I(_02499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05990__A1 (.I(_02499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06085__A4 (.I(_02562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06077__A3 (.I(_02562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06076__A2 (.I(_02562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06073__A2 (.I(_02562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06072__A2 (.I(_02562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06070__A1 (.I(_02562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08549__A2 (.I(_02585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08548__C (.I(_02585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06101__A3 (.I(_02585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06096__A4 (.I(_02585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08755__A1 (.I(_02596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06107__B (.I(_02596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08780__A2 (.I(_02598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08758__A2 (.I(_02598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08750__A3 (.I(_02598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08748__B (.I(_02598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08648__A2 (.I(_02598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06596__A2 (.I(_02598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06119__C (.I(_02598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06110__A2 (.I(_02598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08782__A2 (.I(_02599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06115__B (.I(_02599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06111__B (.I(_02599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08952__A3 (.I(_02604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08926__A2 (.I(_02604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06119__B (.I(_02604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06180__A1 (.I(_02606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06174__A1 (.I(_02606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06168__A1 (.I(_02606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06162__A1 (.I(_02606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06156__A1 (.I(_02606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06150__A1 (.I(_02606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06144__A2 (.I(_02606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06137__A1 (.I(_02606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06126__I (.I(_02606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06125__A3 (.I(_02606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06124__A1 (.I(_02606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06123__A1 (.I(_02606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06688__A1 (.I(_02608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06346__A2 (.I(_02608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06285__A2 (.I(_02608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06284__A2 (.I(_02608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06139__A1 (.I(_02608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06135__A2 (.I(_02608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06124__B1 (.I(_02608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06187__S (.I(_02611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06181__A1 (.I(_02611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06175__A1 (.I(_02611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06169__A1 (.I(_02611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06163__A1 (.I(_02611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06157__A1 (.I(_02611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06151__A1 (.I(_02611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06145__A2 (.I(_02611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06127__A2 (.I(_02611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06196__A3 (.I(_02612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06128__A3 (.I(_02612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09618__A1 (.I(_02619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08890__A1 (.I(_02619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08423__A1 (.I(_02619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07907__A1 (.I(_02619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07570__A1 (.I(_02619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06852__A1 (.I(_02619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06541__A1 (.I(_02619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06245__A1 (.I(_02619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06142__A1 (.I(_02619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08964__A1 (.I(_02621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06138__A1 (.I(_02621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06688__A2 (.I(_02622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06445__A3 (.I(_02622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06368__A3 (.I(_02622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06286__A2 (.I(_02622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06199__A4 (.I(_02622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06138__A2 (.I(_02622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09654__A1 (.I(_02626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09469__A1 (.I(_02626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09451__A1 (.I(_02626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09415__A1 (.I(_02626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09379__A1 (.I(_02626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09318__A1 (.I(_02626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09263__A1 (.I(_02626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09009__A1 (.I(_02626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08984__A1 (.I(_02626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08908__A1 (.I(_02626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07871__A1 (.I(_02626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07833__A1 (.I(_02626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07815__A1 (.I(_02626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06326__A1 (.I(_02626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06227__A1 (.I(_02626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06142__A2 (.I(_02626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06191__A1 (.I(_02628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06190__A2 (.I(_02628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06185__A1 (.I(_02628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06184__A2 (.I(_02628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06179__A1 (.I(_02628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06178__A2 (.I(_02628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06173__A1 (.I(_02628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06172__A2 (.I(_02628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06167__A1 (.I(_02628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06166__A2 (.I(_02628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06161__A1 (.I(_02628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06160__A2 (.I(_02628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06155__A1 (.I(_02628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06154__A2 (.I(_02628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06149__A1 (.I(_02628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06148__A2 (.I(_02628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09317__I (.I(_02631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08983__I (.I(_02631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07943__I (.I(_02631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07606__I (.I(_02631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07274__I (.I(_02631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06906__I (.I(_02631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06540__I (.I(_02631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06192__I (.I(_02631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06147__I (.I(_02631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09364__A1 (.I(_02632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08893__A1 (.I(_02632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08875__A1 (.I(_02632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08026__A1 (.I(_02632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08008__A1 (.I(_02632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07591__A1 (.I(_02632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07375__A1 (.I(_02632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07259__A1 (.I(_02632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07187__A1 (.I(_02632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07169__A1 (.I(_02632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07025__A1 (.I(_02632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06801__A1 (.I(_02632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06569__A1 (.I(_02632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06310__A1 (.I(_02632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06290__A1 (.I(_02632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06149__A2 (.I(_02632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09322__I (.I(_02636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08988__I (.I(_02636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07948__I (.I(_02636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07611__I (.I(_02636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07279__I (.I(_02636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06911__I (.I(_02636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06545__I (.I(_02636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06205__I (.I(_02636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06153__I (.I(_02636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09366__A1 (.I(_02637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08895__A1 (.I(_02637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08877__A1 (.I(_02637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08028__A1 (.I(_02637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08010__A1 (.I(_02637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07593__A1 (.I(_02637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07377__A1 (.I(_02637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07261__A1 (.I(_02637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07189__A1 (.I(_02637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07171__A1 (.I(_02637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07027__A1 (.I(_02637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06803__A1 (.I(_02637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06571__A1 (.I(_02637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06312__A1 (.I(_02637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06292__A1 (.I(_02637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06155__A2 (.I(_02637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09325__I (.I(_02641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08991__I (.I(_02641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07951__I (.I(_02641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07614__I (.I(_02641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07282__I (.I(_02641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06914__I (.I(_02641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06548__I (.I(_02641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06208__I (.I(_02641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06159__I (.I(_02641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09368__A1 (.I(_02642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08897__A1 (.I(_02642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08879__A1 (.I(_02642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08030__A1 (.I(_02642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08012__A1 (.I(_02642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07595__A1 (.I(_02642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07379__A1 (.I(_02642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07263__A1 (.I(_02642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07191__A1 (.I(_02642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07173__A1 (.I(_02642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07029__A1 (.I(_02642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06805__A1 (.I(_02642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06573__A1 (.I(_02642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06314__A1 (.I(_02642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06294__A1 (.I(_02642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06161__A2 (.I(_02642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09328__I (.I(_02646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08994__I (.I(_02646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07954__I (.I(_02646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07617__I (.I(_02646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07285__I (.I(_02646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06917__I (.I(_02646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06551__I (.I(_02646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06211__I (.I(_02646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06165__I (.I(_02646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09370__A1 (.I(_02647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08899__A1 (.I(_02647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08881__A1 (.I(_02647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08032__A1 (.I(_02647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08014__A1 (.I(_02647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07597__A1 (.I(_02647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07381__A1 (.I(_02647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07265__A1 (.I(_02647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07193__A1 (.I(_02647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07175__A1 (.I(_02647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07031__A1 (.I(_02647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06807__A1 (.I(_02647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06575__A1 (.I(_02647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06316__A1 (.I(_02647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06296__A1 (.I(_02647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06167__A2 (.I(_02647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09331__I (.I(_02651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08997__I (.I(_02651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07957__I (.I(_02651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07620__I (.I(_02651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07288__I (.I(_02651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06920__I (.I(_02651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06554__I (.I(_02651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06214__I (.I(_02651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06171__I (.I(_02651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09372__A1 (.I(_02652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08901__A1 (.I(_02652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08883__A1 (.I(_02652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08034__A1 (.I(_02652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08016__A1 (.I(_02652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07599__A1 (.I(_02652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07383__A1 (.I(_02652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07267__A1 (.I(_02652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07195__A1 (.I(_02652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07177__A1 (.I(_02652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07033__A1 (.I(_02652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06809__A1 (.I(_02652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06577__A1 (.I(_02652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06318__A1 (.I(_02652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06298__A1 (.I(_02652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06173__A2 (.I(_02652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09334__I (.I(_02656_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09000__I (.I(_02656_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07960__I (.I(_02656_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07623__I (.I(_02656_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07291__I (.I(_02656_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06923__I (.I(_02656_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06557__I (.I(_02656_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06217__I (.I(_02656_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06177__I (.I(_02656_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09374__A1 (.I(_02657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08903__A1 (.I(_02657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08885__A1 (.I(_02657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08036__A1 (.I(_02657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08018__A1 (.I(_02657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07601__A1 (.I(_02657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07385__A1 (.I(_02657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07269__A1 (.I(_02657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07197__A1 (.I(_02657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07179__A1 (.I(_02657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07035__A1 (.I(_02657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06811__A1 (.I(_02657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06579__A1 (.I(_02657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06320__A1 (.I(_02657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06300__A1 (.I(_02657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06179__A2 (.I(_02657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09337__I (.I(_02661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09003__I (.I(_02661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07963__I (.I(_02661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07626__I (.I(_02661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07294__I (.I(_02661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06926__I (.I(_02661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06560__I (.I(_02661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06220__I (.I(_02661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06183__I (.I(_02661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09376__A1 (.I(_02662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08905__A1 (.I(_02662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08887__A1 (.I(_02662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08038__A1 (.I(_02662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08020__A1 (.I(_02662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07603__A1 (.I(_02662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07387__A1 (.I(_02662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07271__A1 (.I(_02662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07199__A1 (.I(_02662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07181__A1 (.I(_02662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07037__A1 (.I(_02662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06813__A1 (.I(_02662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06581__A1 (.I(_02662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06322__A1 (.I(_02662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06302__A1 (.I(_02662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06185__A2 (.I(_02662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09340__I (.I(_02666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09006__I (.I(_02666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07966__I (.I(_02666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07629__I (.I(_02666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07297__I (.I(_02666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06929__I (.I(_02666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06563__I (.I(_02666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06223__I (.I(_02666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06189__I (.I(_02666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09378__A1 (.I(_02667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08907__A1 (.I(_02667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08889__A1 (.I(_02667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08040__A1 (.I(_02667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08022__A1 (.I(_02667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07605__A1 (.I(_02667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07389__A1 (.I(_02667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07273__A1 (.I(_02667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07201__A1 (.I(_02667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07183__A1 (.I(_02667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07039__A1 (.I(_02667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06815__A1 (.I(_02667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06583__A1 (.I(_02667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06324__A1 (.I(_02667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06304__A1 (.I(_02667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06191__A2 (.I(_02667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09603__A1 (.I(_02669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06525__A1 (.I(_02669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06506__A1 (.I(_02669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06488__A1 (.I(_02669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06469__A1 (.I(_02669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06450__A1 (.I(_02669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06429__A1 (.I(_02669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06410__A1 (.I(_02669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06391__A1 (.I(_02669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06373__A1 (.I(_02669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06351__A1 (.I(_02669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06329__A1 (.I(_02669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06268__A1 (.I(_02669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06248__A1 (.I(_02669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06230__A1 (.I(_02669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06204__A1 (.I(_02669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09379__A2 (.I(_02675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09299__A1 (.I(_02675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09101__A1 (.I(_02675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07925__A1 (.I(_02675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07758__A1 (.I(_02675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07516__A1 (.I(_02675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07130__A1 (.I(_02675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07022__A1 (.I(_02675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06201__A1 (.I(_02675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06200__I (.I(_02676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09672__A1 (.I(_02677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09582__A1 (.I(_02677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09564__A1 (.I(_02677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09546__A1 (.I(_02677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09528__A1 (.I(_02677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09050__A1 (.I(_02677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08762__A1 (.I(_02677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08669__A1 (.I(_02677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07607__A1 (.I(_02677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07004__A1 (.I(_02677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06907__A1 (.I(_02677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06632__A1 (.I(_02677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06614__A1 (.I(_02677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06265__A1 (.I(_02677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06245__A2 (.I(_02677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06201__A2 (.I(_02677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06225__A2 (.I(_02679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06224__A2 (.I(_02679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06222__A2 (.I(_02679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06221__A2 (.I(_02679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06219__A2 (.I(_02679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06218__A2 (.I(_02679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06216__A2 (.I(_02679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06215__A2 (.I(_02679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06213__A2 (.I(_02679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06212__A2 (.I(_02679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06210__A2 (.I(_02679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06209__A2 (.I(_02679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06207__A2 (.I(_02679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06206__A2 (.I(_02679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06204__A2 (.I(_02679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06203__A2 (.I(_02679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09605__A1 (.I(_02681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06527__A1 (.I(_02681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06508__A1 (.I(_02681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06490__A1 (.I(_02681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06471__A1 (.I(_02681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06452__A1 (.I(_02681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06431__A1 (.I(_02681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06412__A1 (.I(_02681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06393__A1 (.I(_02681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06375__A1 (.I(_02681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06353__A1 (.I(_02681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06331__A1 (.I(_02681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06270__A1 (.I(_02681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06250__A1 (.I(_02681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06232__A1 (.I(_02681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06207__A1 (.I(_02681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09607__A1 (.I(_02683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06529__A1 (.I(_02683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06510__A1 (.I(_02683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06492__A1 (.I(_02683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06473__A1 (.I(_02683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06454__A1 (.I(_02683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06433__A1 (.I(_02683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06414__A1 (.I(_02683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06395__A1 (.I(_02683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06377__A1 (.I(_02683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06355__A1 (.I(_02683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06333__A1 (.I(_02683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06272__A1 (.I(_02683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06252__A1 (.I(_02683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06234__A1 (.I(_02683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06210__A1 (.I(_02683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09609__A1 (.I(_02685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06531__A1 (.I(_02685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06512__A1 (.I(_02685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06494__A1 (.I(_02685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06475__A1 (.I(_02685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06456__A1 (.I(_02685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06435__A1 (.I(_02685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06416__A1 (.I(_02685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06397__A1 (.I(_02685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06379__A1 (.I(_02685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06357__A1 (.I(_02685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06335__A1 (.I(_02685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06274__A1 (.I(_02685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06254__A1 (.I(_02685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06236__A1 (.I(_02685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06213__A1 (.I(_02685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09611__A1 (.I(_02687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06533__A1 (.I(_02687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06514__A1 (.I(_02687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06496__A1 (.I(_02687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06477__A1 (.I(_02687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06458__A1 (.I(_02687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06437__A1 (.I(_02687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06418__A1 (.I(_02687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06399__A1 (.I(_02687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06381__A1 (.I(_02687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06359__A1 (.I(_02687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06337__A1 (.I(_02687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06276__A1 (.I(_02687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06256__A1 (.I(_02687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06238__A1 (.I(_02687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06216__A1 (.I(_02687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09613__A1 (.I(_02689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06535__A1 (.I(_02689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06516__A1 (.I(_02689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06498__A1 (.I(_02689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06479__A1 (.I(_02689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06460__A1 (.I(_02689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06439__A1 (.I(_02689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06420__A1 (.I(_02689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06401__A1 (.I(_02689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06383__A1 (.I(_02689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06361__A1 (.I(_02689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06339__A1 (.I(_02689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06278__A1 (.I(_02689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06258__A1 (.I(_02689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06240__A1 (.I(_02689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06219__A1 (.I(_02689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09615__A1 (.I(_02691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06537__A1 (.I(_02691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06518__A1 (.I(_02691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06500__A1 (.I(_02691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06481__A1 (.I(_02691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06462__A1 (.I(_02691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06441__A1 (.I(_02691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06422__A1 (.I(_02691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06403__A1 (.I(_02691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06385__A1 (.I(_02691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06363__A1 (.I(_02691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06341__A1 (.I(_02691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06280__A1 (.I(_02691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06260__A1 (.I(_02691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06242__A1 (.I(_02691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06222__A1 (.I(_02691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09617__A1 (.I(_02693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06539__A1 (.I(_02693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06520__A1 (.I(_02693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06502__A1 (.I(_02693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06483__A1 (.I(_02693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06464__A1 (.I(_02693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06443__A1 (.I(_02693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06424__A1 (.I(_02693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06405__A1 (.I(_02693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06387__A1 (.I(_02693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06365__A1 (.I(_02693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06343__A1 (.I(_02693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06282__A1 (.I(_02693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06262__A1 (.I(_02693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06244__A1 (.I(_02693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06225__A1 (.I(_02693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08965__A1 (.I(_02695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08248__A1 (.I(_02695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08113__A1 (.I(_02695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07444__A1 (.I(_02695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06870__A1 (.I(_02695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06689__A1 (.I(_02695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06632__A2 (.I(_02695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06287__A1 (.I(_02695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06227__A2 (.I(_02695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06244__A2 (.I(_02697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06243__A2 (.I(_02697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06242__A2 (.I(_02697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06241__A2 (.I(_02697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06240__A2 (.I(_02697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06239__A2 (.I(_02697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06238__A2 (.I(_02697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06237__A2 (.I(_02697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06236__A2 (.I(_02697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06235__A2 (.I(_02697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06234__A2 (.I(_02697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06233__A2 (.I(_02697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06232__A2 (.I(_02697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06231__A2 (.I(_02697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06230__A2 (.I(_02697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06229__A2 (.I(_02697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06262__A2 (.I(_02707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06261__A2 (.I(_02707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06260__A2 (.I(_02707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06259__A2 (.I(_02707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06258__A2 (.I(_02707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06257__A2 (.I(_02707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06256__A2 (.I(_02707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06255__A2 (.I(_02707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06254__A2 (.I(_02707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06253__A2 (.I(_02707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06252__A2 (.I(_02707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06251__A2 (.I(_02707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06250__A2 (.I(_02707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06249__A2 (.I(_02707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06248__A2 (.I(_02707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06247__A2 (.I(_02707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09636__A1 (.I(_02717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09318__A2 (.I(_02717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08095__A1 (.I(_02717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07776__A1 (.I(_02717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07534__A1 (.I(_02717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07148__A1 (.I(_02717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06816__A1 (.I(_02717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06566__A1 (.I(_02717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06265__A2 (.I(_02717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06282__A2 (.I(_02719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06281__A2 (.I(_02719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06280__A2 (.I(_02719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06279__A2 (.I(_02719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06278__A2 (.I(_02719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06277__A2 (.I(_02719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06276__A2 (.I(_02719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06275__A2 (.I(_02719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06274__A2 (.I(_02719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06273__A2 (.I(_02719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06272__A2 (.I(_02719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06271__A2 (.I(_02719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06270__A2 (.I(_02719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06269__A2 (.I(_02719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06268__A2 (.I(_02719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06267__A2 (.I(_02719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08949__A1 (.I(_02728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08938__A1 (.I(_02728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06669__A1 (.I(_02728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06445__A1 (.I(_02728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06346__A1 (.I(_02728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06285__A1 (.I(_02728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09600__A1 (.I(_02731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09361__A1 (.I(_02731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08890__A2 (.I(_02731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08872__A1 (.I(_02731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08023__A1 (.I(_02731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08005__A1 (.I(_02731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07588__A1 (.I(_02731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07372__A1 (.I(_02731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07256__A1 (.I(_02731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07184__A1 (.I(_02731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07166__A1 (.I(_02731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07022__A2 (.I(_02731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06798__A1 (.I(_02731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06566__A2 (.I(_02731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06307__A1 (.I(_02731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06287__A2 (.I(_02731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06304__A2 (.I(_02733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06303__A2 (.I(_02733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06302__A2 (.I(_02733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06301__A2 (.I(_02733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06300__A2 (.I(_02733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06299__A2 (.I(_02733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06298__A2 (.I(_02733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06297__A2 (.I(_02733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06296__A2 (.I(_02733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06295__A2 (.I(_02733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06294__A2 (.I(_02733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06293__A2 (.I(_02733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06292__A2 (.I(_02733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06291__A2 (.I(_02733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06290__A2 (.I(_02733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06289__A2 (.I(_02733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09672__A2 (.I(_02743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09451__A2 (.I(_02743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09137__A1 (.I(_02743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07480__A1 (.I(_02743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07408__A1 (.I(_02743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07318__A1 (.I(_02743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07094__A1 (.I(_02743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06670__A1 (.I(_02743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06307__A2 (.I(_02743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06324__A2 (.I(_02745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06323__A2 (.I(_02745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06322__A2 (.I(_02745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06321__A2 (.I(_02745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06320__A2 (.I(_02745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06319__A2 (.I(_02745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06318__A2 (.I(_02745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06317__A2 (.I(_02745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06316__A2 (.I(_02745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06315__A2 (.I(_02745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06314__A2 (.I(_02745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06313__A2 (.I(_02745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06312__A2 (.I(_02745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06311__A2 (.I(_02745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06310__A2 (.I(_02745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06309__A2 (.I(_02745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09600__A2 (.I(_02754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09027__A1 (.I(_02754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08651__A1 (.I(_02754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08041__A1 (.I(_02754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07632__A1 (.I(_02754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06888__A1 (.I(_02754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06614__A2 (.I(_02754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06503__A1 (.I(_02754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06326__A2 (.I(_02754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06343__A2 (.I(_02756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06342__A2 (.I(_02756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06341__A2 (.I(_02756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06340__A2 (.I(_02756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06339__A2 (.I(_02756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06338__A2 (.I(_02756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06337__A2 (.I(_02756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06336__A2 (.I(_02756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06335__A2 (.I(_02756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06334__A2 (.I(_02756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06333__A2 (.I(_02756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06332__A2 (.I(_02756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06331__A2 (.I(_02756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06330__A2 (.I(_02756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06329__A2 (.I(_02756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06328__A2 (.I(_02756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09397__A1 (.I(_02766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08984__A2 (.I(_02766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08762__A2 (.I(_02766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07668__A1 (.I(_02766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07372__A2 (.I(_02766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07202__A1 (.I(_02766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06950__A1 (.I(_02766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06388__A1 (.I(_02766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06348__A1 (.I(_02766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06347__I (.I(_02767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09299__A2 (.I(_02768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09191__A1 (.I(_02768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07336__A1 (.I(_02768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07318__A2 (.I(_02768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07300__A1 (.I(_02768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07275__A1 (.I(_02768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06888__A2 (.I(_02768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06870__A2 (.I(_02768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06852__A2 (.I(_02768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06834__A1 (.I(_02768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06816__A2 (.I(_02768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06779__A1 (.I(_02768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06761__A1 (.I(_02768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06743__A1 (.I(_02768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06725__A1 (.I(_02768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06348__A2 (.I(_02768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06365__A2 (.I(_02770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06364__A2 (.I(_02770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06363__A2 (.I(_02770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06362__A2 (.I(_02770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06361__A2 (.I(_02770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06360__A2 (.I(_02770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06359__A2 (.I(_02770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06358__A2 (.I(_02770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06357__A2 (.I(_02770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06356__A2 (.I(_02770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06355__A2 (.I(_02770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06354__A2 (.I(_02770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06353__A2 (.I(_02770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06352__A2 (.I(_02770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06351__A2 (.I(_02770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06350__A2 (.I(_02770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09546__A2 (.I(_02780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09361__A2 (.I(_02780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09227__A1 (.I(_02780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08059__A1 (.I(_02780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07833__A2 (.I(_02780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07390__A1 (.I(_02780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07040__A1 (.I(_02780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06743__A2 (.I(_02780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06370__A1 (.I(_02780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08651__A2 (.I(_02782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08113__A2 (.I(_02782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07907__A2 (.I(_02782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07889__A1 (.I(_02782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07776__A2 (.I(_02782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07758__A2 (.I(_02782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07740__A1 (.I(_02782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07408__A2 (.I(_02782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06651__A1 (.I(_02782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06522__A1 (.I(_02782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06485__A1 (.I(_02782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06466__A1 (.I(_02782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06426__A1 (.I(_02782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06407__A1 (.I(_02782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06388__A2 (.I(_02782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06370__A2 (.I(_02782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06387__A2 (.I(_02784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06386__A2 (.I(_02784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06385__A2 (.I(_02784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06384__A2 (.I(_02784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06383__A2 (.I(_02784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06382__A2 (.I(_02784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06381__A2 (.I(_02784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06380__A2 (.I(_02784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06379__A2 (.I(_02784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06378__A2 (.I(_02784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06377__A2 (.I(_02784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06376__A2 (.I(_02784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06375__A2 (.I(_02784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06374__A2 (.I(_02784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06373__A2 (.I(_02784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06372__A2 (.I(_02784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06405__A2 (.I(_02794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06404__A2 (.I(_02794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06403__A2 (.I(_02794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06402__A2 (.I(_02794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06401__A2 (.I(_02794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06400__A2 (.I(_02794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06399__A2 (.I(_02794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06398__A2 (.I(_02794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06397__A2 (.I(_02794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06396__A2 (.I(_02794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06395__A2 (.I(_02794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06394__A2 (.I(_02794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06393__A2 (.I(_02794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06392__A2 (.I(_02794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06391__A2 (.I(_02794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06390__A2 (.I(_02794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08908__A2 (.I(_02803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08854__A1 (.I(_02803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07686__A1 (.I(_02803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07256__A2 (.I(_02803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07220__A1 (.I(_02803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06968__A1 (.I(_02803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06907__A2 (.I(_02803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06725__A2 (.I(_02803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06407__A2 (.I(_02803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06424__A2 (.I(_02805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06423__A2 (.I(_02805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06422__A2 (.I(_02805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06421__A2 (.I(_02805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06420__A2 (.I(_02805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06419__A2 (.I(_02805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06418__A2 (.I(_02805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06417__A2 (.I(_02805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06416__A2 (.I(_02805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06415__A2 (.I(_02805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06414__A2 (.I(_02805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06413__A2 (.I(_02805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06412__A2 (.I(_02805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06411__A2 (.I(_02805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06410__A2 (.I(_02805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06409__A2 (.I(_02805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09281__A1 (.I(_02814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09050__A2 (.I(_02814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07871__A2 (.I(_02814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07704__A1 (.I(_02814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07588__A2 (.I(_02814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07238__A1 (.I(_02814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06986__A1 (.I(_02814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06761__A2 (.I(_02814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06426__A2 (.I(_02814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06443__A2 (.I(_02816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06442__A2 (.I(_02816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06441__A2 (.I(_02816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06440__A2 (.I(_02816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06439__A2 (.I(_02816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06438__A2 (.I(_02816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06437__A2 (.I(_02816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06436__A2 (.I(_02816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06435__A2 (.I(_02816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06434__A2 (.I(_02816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06433__A2 (.I(_02816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06432__A2 (.I(_02816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06431__A2 (.I(_02816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06430__A2 (.I(_02816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06429__A2 (.I(_02816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06428__A2 (.I(_02816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09263__A2 (.I(_02825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09173__A1 (.I(_02825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08872__A2 (.I(_02825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08077__A1 (.I(_02825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07889__A2 (.I(_02825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07552__A1 (.I(_02825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07004__A2 (.I(_02825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06834__A2 (.I(_02825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06447__A1 (.I(_02825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09343__A1 (.I(_02827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07444__A2 (.I(_02827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07148__A2 (.I(_02827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07130__A2 (.I(_02827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07112__A1 (.I(_02827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07094__A2 (.I(_02827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07076__A1 (.I(_02827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07058__A1 (.I(_02827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07040__A2 (.I(_02827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06986__A2 (.I(_02827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06968__A2 (.I(_02827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06950__A2 (.I(_02827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06932__A1 (.I(_02827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06541__A2 (.I(_02827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06503__A2 (.I(_02827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06447__A2 (.I(_02827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06464__A2 (.I(_02829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06463__A2 (.I(_02829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06462__A2 (.I(_02829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06461__A2 (.I(_02829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06460__A2 (.I(_02829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06459__A2 (.I(_02829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06458__A2 (.I(_02829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06457__A2 (.I(_02829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06456__A2 (.I(_02829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06455__A2 (.I(_02829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06454__A2 (.I(_02829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06453__A2 (.I(_02829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06452__A2 (.I(_02829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06451__A2 (.I(_02829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06450__A2 (.I(_02829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06449__A2 (.I(_02829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09654__A2 (.I(_02838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09564__A2 (.I(_02838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09209__A1 (.I(_02838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07987__A1 (.I(_02838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07426__A1 (.I(_02838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07300__A2 (.I(_02838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07166__A2 (.I(_02838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07058__A2 (.I(_02838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06466__A2 (.I(_02838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06483__A2 (.I(_02840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06482__A2 (.I(_02840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06481__A2 (.I(_02840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06480__A2 (.I(_02840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06479__A2 (.I(_02840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06478__A2 (.I(_02840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06477__A2 (.I(_02840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06476__A2 (.I(_02840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06475__A2 (.I(_02840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06474__A2 (.I(_02840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06473__A2 (.I(_02840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06472__A2 (.I(_02840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06471__A2 (.I(_02840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06470__A2 (.I(_02840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06469__A2 (.I(_02840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06468__A2 (.I(_02840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09528__A2 (.I(_02849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09343__A2 (.I(_02849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09245__A1 (.I(_02849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08023__A2 (.I(_02849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07815__A2 (.I(_02849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07722__A1 (.I(_02849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06779__A2 (.I(_02849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06707__A1 (.I(_02849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06485__A2 (.I(_02849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06502__A2 (.I(_02851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06501__A2 (.I(_02851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06500__A2 (.I(_02851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06499__A2 (.I(_02851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06498__A2 (.I(_02851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06497__A2 (.I(_02851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06496__A2 (.I(_02851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06495__A2 (.I(_02851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06494__A2 (.I(_02851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06493__A2 (.I(_02851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06492__A2 (.I(_02851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06491__A2 (.I(_02851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06490__A2 (.I(_02851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06489__A2 (.I(_02851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06488__A2 (.I(_02851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06487__A2 (.I(_02851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06520__A2 (.I(_02861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06519__A2 (.I(_02861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06518__A2 (.I(_02861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06517__A2 (.I(_02861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06516__A2 (.I(_02861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06515__A2 (.I(_02861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06514__A2 (.I(_02861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06513__A2 (.I(_02861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06512__A2 (.I(_02861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06511__A2 (.I(_02861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06510__A2 (.I(_02861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06509__A2 (.I(_02861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06508__A2 (.I(_02861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06507__A2 (.I(_02861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06506__A2 (.I(_02861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06505__A2 (.I(_02861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09433__A1 (.I(_02870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09191__A2 (.I(_02870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09009__A2 (.I(_02870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08669__A2 (.I(_02870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07650__A1 (.I(_02870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07354__A1 (.I(_02870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07184__A2 (.I(_02870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06932__A2 (.I(_02870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06522__A2 (.I(_02870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06539__A2 (.I(_02872_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06538__A2 (.I(_02872_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06537__A2 (.I(_02872_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06536__A2 (.I(_02872_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06535__A2 (.I(_02872_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06534__A2 (.I(_02872_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06533__A2 (.I(_02872_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06532__A2 (.I(_02872_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06531__A2 (.I(_02872_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06530__A2 (.I(_02872_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06529__A2 (.I(_02872_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06528__A2 (.I(_02872_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06527__A2 (.I(_02872_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06526__A2 (.I(_02872_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06525__A2 (.I(_02872_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06524__A2 (.I(_02872_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06891__A1 (.I(_02881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06873__A1 (.I(_02881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06855__A1 (.I(_02881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06837__A1 (.I(_02881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06819__A1 (.I(_02881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06782__A1 (.I(_02881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06764__A1 (.I(_02881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06746__A1 (.I(_02881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06728__A1 (.I(_02881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06710__A1 (.I(_02881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06692__A1 (.I(_02881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06673__A1 (.I(_02881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06654__A1 (.I(_02881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06635__A1 (.I(_02881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06617__A1 (.I(_02881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06544__A1 (.I(_02881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06565__A2 (.I(_02883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06564__A2 (.I(_02883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06562__A2 (.I(_02883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06561__A2 (.I(_02883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06559__A2 (.I(_02883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06558__A2 (.I(_02883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06556__A2 (.I(_02883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06555__A2 (.I(_02883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06553__A2 (.I(_02883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06552__A2 (.I(_02883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06550__A2 (.I(_02883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06549__A2 (.I(_02883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06547__A2 (.I(_02883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06546__A2 (.I(_02883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06544__A2 (.I(_02883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06543__A2 (.I(_02883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06893__A1 (.I(_02885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06875__A1 (.I(_02885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06857__A1 (.I(_02885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06839__A1 (.I(_02885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06821__A1 (.I(_02885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06784__A1 (.I(_02885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06766__A1 (.I(_02885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06748__A1 (.I(_02885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06730__A1 (.I(_02885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06712__A1 (.I(_02885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06694__A1 (.I(_02885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06675__A1 (.I(_02885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06656__A1 (.I(_02885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06637__A1 (.I(_02885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06619__A1 (.I(_02885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06547__A1 (.I(_02885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06895__A1 (.I(_02887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06877__A1 (.I(_02887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06859__A1 (.I(_02887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06841__A1 (.I(_02887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06823__A1 (.I(_02887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06786__A1 (.I(_02887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06768__A1 (.I(_02887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06750__A1 (.I(_02887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06732__A1 (.I(_02887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06714__A1 (.I(_02887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06696__A1 (.I(_02887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06677__A1 (.I(_02887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06658__A1 (.I(_02887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06639__A1 (.I(_02887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06621__A1 (.I(_02887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06550__A1 (.I(_02887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06897__A1 (.I(_02889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06879__A1 (.I(_02889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06861__A1 (.I(_02889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06843__A1 (.I(_02889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06825__A1 (.I(_02889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06788__A1 (.I(_02889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06770__A1 (.I(_02889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06752__A1 (.I(_02889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06734__A1 (.I(_02889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06716__A1 (.I(_02889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06698__A1 (.I(_02889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06679__A1 (.I(_02889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06660__A1 (.I(_02889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06641__A1 (.I(_02889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06623__A1 (.I(_02889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06553__A1 (.I(_02889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06899__A1 (.I(_02891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06881__A1 (.I(_02891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06863__A1 (.I(_02891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06845__A1 (.I(_02891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06827__A1 (.I(_02891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06790__A1 (.I(_02891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06772__A1 (.I(_02891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06754__A1 (.I(_02891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06736__A1 (.I(_02891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06718__A1 (.I(_02891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06700__A1 (.I(_02891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06681__A1 (.I(_02891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06662__A1 (.I(_02891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06643__A1 (.I(_02891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06625__A1 (.I(_02891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06556__A1 (.I(_02891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06901__A1 (.I(_02893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06883__A1 (.I(_02893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06865__A1 (.I(_02893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06847__A1 (.I(_02893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06829__A1 (.I(_02893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06792__A1 (.I(_02893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06774__A1 (.I(_02893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06756__A1 (.I(_02893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06738__A1 (.I(_02893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06720__A1 (.I(_02893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06702__A1 (.I(_02893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06683__A1 (.I(_02893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06664__A1 (.I(_02893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06645__A1 (.I(_02893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06627__A1 (.I(_02893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06559__A1 (.I(_02893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06903__A1 (.I(_02895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06885__A1 (.I(_02895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06867__A1 (.I(_02895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06849__A1 (.I(_02895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06831__A1 (.I(_02895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06794__A1 (.I(_02895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06776__A1 (.I(_02895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06758__A1 (.I(_02895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06740__A1 (.I(_02895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06722__A1 (.I(_02895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06704__A1 (.I(_02895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06685__A1 (.I(_02895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06666__A1 (.I(_02895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06647__A1 (.I(_02895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06629__A1 (.I(_02895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06562__A1 (.I(_02895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06905__A1 (.I(_02897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06887__A1 (.I(_02897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06869__A1 (.I(_02897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06851__A1 (.I(_02897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06833__A1 (.I(_02897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06796__A1 (.I(_02897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06778__A1 (.I(_02897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06760__A1 (.I(_02897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06742__A1 (.I(_02897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06724__A1 (.I(_02897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06706__A1 (.I(_02897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06687__A1 (.I(_02897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06668__A1 (.I(_02897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06649__A1 (.I(_02897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06631__A1 (.I(_02897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06565__A1 (.I(_02897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06583__A2 (.I(_02900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06582__A2 (.I(_02900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06581__A2 (.I(_02900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06580__A2 (.I(_02900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06579__A2 (.I(_02900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06578__A2 (.I(_02900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06577__A2 (.I(_02900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06576__A2 (.I(_02900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06575__A2 (.I(_02900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06574__A2 (.I(_02900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06573__A2 (.I(_02900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06572__A2 (.I(_02900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06571__A2 (.I(_02900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06570__A2 (.I(_02900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06569__A2 (.I(_02900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06568__A2 (.I(_02900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08612__A1 (.I(_02909_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08611__A1 (.I(_02909_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08374__A1 (.I(_02909_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08355__A1 (.I(_02909_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08349__A1 (.I(_02909_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08332__A1 (.I(_02909_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08307__A1 (.I(_02909_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08300__A1 (.I(_02909_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08289__A1 (.I(_02909_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08286__A1 (.I(_02909_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08280__A1 (.I(_02909_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08266__A1 (.I(_02909_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06586__A1 (.I(_02909_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09099__S (.I(_02910_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09068__I (.I(_02910_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06586__B (.I(_02910_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08568__B (.I(_02911_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08397__A1 (.I(_02911_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08340__A1 (.I(_02911_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08333__A1 (.I(_02911_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08329__I (.I(_02911_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06587__B (.I(_02911_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09700__A1 (.I(_02912_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06610__A1 (.I(_02912_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06604__A1 (.I(_02912_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06588__A2 (.I(_02912_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08755__A2 (.I(_02914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08754__C (.I(_02914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07794__A2 (.I(_02914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06591__A2 (.I(_02914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08166__A2 (.I(_02915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08163__A1 (.I(_02915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08159__A1 (.I(_02915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08158__A2 (.I(_02915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08151__B (.I(_02915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08150__A2 (.I(_02915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08144__B (.I(_02915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08143__A2 (.I(_02915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08137__A2 (.I(_02915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08135__A2 (.I(_02915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06595__A1 (.I(_02915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06597__A2 (.I(_02920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08171__B2 (.I(_02922_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06599__A3 (.I(_02922_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08246__A2 (.I(_02924_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08244__A2 (.I(_02924_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08234__A2 (.I(_02924_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08231__A1 (.I(_02924_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08164__A1 (.I(_02924_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08155__A2 (.I(_02924_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08154__B (.I(_02924_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08148__A2 (.I(_02924_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08147__B (.I(_02924_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08137__B (.I(_02924_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06601__B (.I(_02924_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09701__A1 (.I(_02927_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07806__A2 (.I(_02927_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06610__A2 (.I(_02927_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06604__A2 (.I(_02927_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06609__A2 (.I(_02929_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06608__A2 (.I(_02929_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06607__A3 (.I(_02929_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06631__A2 (.I(_02935_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06630__A2 (.I(_02935_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06629__A2 (.I(_02935_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06628__A2 (.I(_02935_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06627__A2 (.I(_02935_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06626__A2 (.I(_02935_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06625__A2 (.I(_02935_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06624__A2 (.I(_02935_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06623__A2 (.I(_02935_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06622__A2 (.I(_02935_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06621__A2 (.I(_02935_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06620__A2 (.I(_02935_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06619__A2 (.I(_02935_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06618__A2 (.I(_02935_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06617__A2 (.I(_02935_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06616__A2 (.I(_02935_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06649__A2 (.I(_02945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06648__A2 (.I(_02945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06647__A2 (.I(_02945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06646__A2 (.I(_02945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06645__A2 (.I(_02945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06644__A2 (.I(_02945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06643__A2 (.I(_02945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06642__A2 (.I(_02945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06641__A2 (.I(_02945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06640__A2 (.I(_02945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06639__A2 (.I(_02945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06638__A2 (.I(_02945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06637__A2 (.I(_02945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06636__A2 (.I(_02945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06635__A2 (.I(_02945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06634__A2 (.I(_02945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09582__A2 (.I(_02954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09469__A2 (.I(_02954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09155__A1 (.I(_02954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08005__A2 (.I(_02954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07944__A1 (.I(_02954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07462__A1 (.I(_02954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07275__A2 (.I(_02954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07076__A2 (.I(_02954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06651__A2 (.I(_02954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06668__A2 (.I(_02956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06667__A2 (.I(_02956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06666__A2 (.I(_02956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06665__A2 (.I(_02956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06664__A2 (.I(_02956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06663__A2 (.I(_02956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06662__A2 (.I(_02956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06661__A2 (.I(_02956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06660__A2 (.I(_02956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06659__A2 (.I(_02956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06658__A2 (.I(_02956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06657__A2 (.I(_02956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06656__A2 (.I(_02956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06655__A2 (.I(_02956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06654__A2 (.I(_02956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06653__A2 (.I(_02956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08423__A2 (.I(_02965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08248__A2 (.I(_02965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08095__A2 (.I(_02965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08077__A2 (.I(_02965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08059__A2 (.I(_02965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08041__A2 (.I(_02965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07987__A2 (.I(_02965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07969__A1 (.I(_02965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07944__A2 (.I(_02965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07925__A2 (.I(_02965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07722__A2 (.I(_02965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07704__A2 (.I(_02965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07686__A2 (.I(_02965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07668__A2 (.I(_02965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07650__A2 (.I(_02965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06670__A2 (.I(_02965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06687__A2 (.I(_02967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06686__A2 (.I(_02967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06685__A2 (.I(_02967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06684__A2 (.I(_02967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06683__A2 (.I(_02967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06682__A2 (.I(_02967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06681__A2 (.I(_02967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06680__A2 (.I(_02967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06679__A2 (.I(_02967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06678__A2 (.I(_02967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06677__A2 (.I(_02967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06676__A2 (.I(_02967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06675__A2 (.I(_02967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06674__A2 (.I(_02967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06673__A2 (.I(_02967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06672__A2 (.I(_02967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07632__A2 (.I(_02976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07570__A2 (.I(_02976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07552__A2 (.I(_02976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07534__A2 (.I(_02976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07516__A2 (.I(_02976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07498__A1 (.I(_02976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07480__A2 (.I(_02976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07462__A2 (.I(_02976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07426__A2 (.I(_02976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07390__A2 (.I(_02976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07354__A2 (.I(_02976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07238__A2 (.I(_02976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07220__A2 (.I(_02976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07202__A2 (.I(_02976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06707__A2 (.I(_02976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06689__A2 (.I(_02976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06706__A2 (.I(_02978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06705__A2 (.I(_02978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06704__A2 (.I(_02978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06703__A2 (.I(_02978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06702__A2 (.I(_02978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06701__A2 (.I(_02978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06700__A2 (.I(_02978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06699__A2 (.I(_02978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06698__A2 (.I(_02978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06697__A2 (.I(_02978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06696__A2 (.I(_02978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06695__A2 (.I(_02978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06694__A2 (.I(_02978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06693__A2 (.I(_02978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06692__A2 (.I(_02978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06691__A2 (.I(_02978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06724__A2 (.I(_02988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06723__A2 (.I(_02988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06722__A2 (.I(_02988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06721__A2 (.I(_02988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06720__A2 (.I(_02988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06719__A2 (.I(_02988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06718__A2 (.I(_02988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06717__A2 (.I(_02988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06716__A2 (.I(_02988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06715__A2 (.I(_02988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06714__A2 (.I(_02988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06713__A2 (.I(_02988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06712__A2 (.I(_02988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06711__A2 (.I(_02988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06710__A2 (.I(_02988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06709__A2 (.I(_02988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06742__A2 (.I(_02998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06741__A2 (.I(_02998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06740__A2 (.I(_02998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06739__A2 (.I(_02998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06738__A2 (.I(_02998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06737__A2 (.I(_02998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06736__A2 (.I(_02998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06735__A2 (.I(_02998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06734__A2 (.I(_02998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06733__A2 (.I(_02998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06732__A2 (.I(_02998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06731__A2 (.I(_02998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06730__A2 (.I(_02998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06729__A2 (.I(_02998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06728__A2 (.I(_02998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06727__A2 (.I(_02998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06760__A2 (.I(_03008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06759__A2 (.I(_03008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06758__A2 (.I(_03008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06757__A2 (.I(_03008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06756__A2 (.I(_03008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06755__A2 (.I(_03008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06754__A2 (.I(_03008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06753__A2 (.I(_03008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06752__A2 (.I(_03008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06751__A2 (.I(_03008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06750__A2 (.I(_03008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06749__A2 (.I(_03008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06748__A2 (.I(_03008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06747__A2 (.I(_03008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06746__A2 (.I(_03008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06745__A2 (.I(_03008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06778__A2 (.I(_03018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06777__A2 (.I(_03018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06776__A2 (.I(_03018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06775__A2 (.I(_03018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06774__A2 (.I(_03018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06773__A2 (.I(_03018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06772__A2 (.I(_03018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06771__A2 (.I(_03018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06770__A2 (.I(_03018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06769__A2 (.I(_03018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06768__A2 (.I(_03018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06767__A2 (.I(_03018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06766__A2 (.I(_03018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06765__A2 (.I(_03018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06764__A2 (.I(_03018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06763__A2 (.I(_03018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06796__A2 (.I(_03028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06795__A2 (.I(_03028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06794__A2 (.I(_03028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06793__A2 (.I(_03028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06792__A2 (.I(_03028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06791__A2 (.I(_03028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06790__A2 (.I(_03028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06789__A2 (.I(_03028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06788__A2 (.I(_03028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06787__A2 (.I(_03028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06786__A2 (.I(_03028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06785__A2 (.I(_03028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06784__A2 (.I(_03028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06783__A2 (.I(_03028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06782__A2 (.I(_03028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06781__A2 (.I(_03028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09415__A2 (.I(_03037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09119__A1 (.I(_03037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07969__A2 (.I(_03037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07740__A2 (.I(_03037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07607__A2 (.I(_03037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07498__A2 (.I(_03037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07336__A2 (.I(_03037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07112__A2 (.I(_03037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06798__A2 (.I(_03037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06815__A2 (.I(_03039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06814__A2 (.I(_03039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06813__A2 (.I(_03039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06812__A2 (.I(_03039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06811__A2 (.I(_03039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06810__A2 (.I(_03039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06809__A2 (.I(_03039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06808__A2 (.I(_03039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06807__A2 (.I(_03039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06806__A2 (.I(_03039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06805__A2 (.I(_03039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06804__A2 (.I(_03039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06803__A2 (.I(_03039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06802__A2 (.I(_03039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06801__A2 (.I(_03039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06800__A2 (.I(_03039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06833__A2 (.I(_03049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06832__A2 (.I(_03049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06831__A2 (.I(_03049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06830__A2 (.I(_03049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06829__A2 (.I(_03049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06828__A2 (.I(_03049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06827__A2 (.I(_03049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06826__A2 (.I(_03049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06825__A2 (.I(_03049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06824__A2 (.I(_03049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06823__A2 (.I(_03049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06822__A2 (.I(_03049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06821__A2 (.I(_03049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06820__A2 (.I(_03049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06819__A2 (.I(_03049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06818__A2 (.I(_03049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06835__I (.I(_03058_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06851__A2 (.I(_03059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06850__A2 (.I(_03059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06849__A2 (.I(_03059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06848__A2 (.I(_03059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06847__A2 (.I(_03059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06846__A2 (.I(_03059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06845__A2 (.I(_03059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06844__A2 (.I(_03059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06843__A2 (.I(_03059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06842__A2 (.I(_03059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06841__A2 (.I(_03059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06840__A2 (.I(_03059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06839__A2 (.I(_03059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06838__A2 (.I(_03059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06837__A2 (.I(_03059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06836__A2 (.I(_03059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06853__I (.I(_03068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06869__A2 (.I(_03069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06868__A2 (.I(_03069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06867__A2 (.I(_03069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06866__A2 (.I(_03069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06865__A2 (.I(_03069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06864__A2 (.I(_03069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06863__A2 (.I(_03069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06862__A2 (.I(_03069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06861__A2 (.I(_03069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06860__A2 (.I(_03069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06859__A2 (.I(_03069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06858__A2 (.I(_03069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06857__A2 (.I(_03069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06856__A2 (.I(_03069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06855__A2 (.I(_03069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06854__A2 (.I(_03069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06887__A2 (.I(_03079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06886__A2 (.I(_03079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06885__A2 (.I(_03079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06884__A2 (.I(_03079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06883__A2 (.I(_03079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06882__A2 (.I(_03079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06881__A2 (.I(_03079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06880__A2 (.I(_03079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06879__A2 (.I(_03079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06878__A2 (.I(_03079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06877__A2 (.I(_03079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06876__A2 (.I(_03079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06875__A2 (.I(_03079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06874__A2 (.I(_03079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06873__A2 (.I(_03079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06872__A2 (.I(_03079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06905__A2 (.I(_03089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06904__A2 (.I(_03089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06903__A2 (.I(_03089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06902__A2 (.I(_03089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06901__A2 (.I(_03089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06900__A2 (.I(_03089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06899__A2 (.I(_03089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06898__A2 (.I(_03089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06897__A2 (.I(_03089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06896__A2 (.I(_03089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06895__A2 (.I(_03089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06894__A2 (.I(_03089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06893__A2 (.I(_03089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06892__A2 (.I(_03089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06891__A2 (.I(_03089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06890__A2 (.I(_03089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07241__A1 (.I(_03098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07223__A1 (.I(_03098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07205__A1 (.I(_03098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07151__A1 (.I(_03098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07133__A1 (.I(_03098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07115__A1 (.I(_03098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07097__A1 (.I(_03098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07079__A1 (.I(_03098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07061__A1 (.I(_03098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07043__A1 (.I(_03098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07007__A1 (.I(_03098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06989__A1 (.I(_03098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06971__A1 (.I(_03098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06953__A1 (.I(_03098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06935__A1 (.I(_03098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06910__A1 (.I(_03098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06931__A2 (.I(_03100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06930__A2 (.I(_03100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06928__A2 (.I(_03100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06927__A2 (.I(_03100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06925__A2 (.I(_03100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06924__A2 (.I(_03100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06922__A2 (.I(_03100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06921__A2 (.I(_03100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06919__A2 (.I(_03100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06918__A2 (.I(_03100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06916__A2 (.I(_03100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06915__A2 (.I(_03100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06913__A2 (.I(_03100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06912__A2 (.I(_03100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06910__A2 (.I(_03100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06909__A2 (.I(_03100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07243__A1 (.I(_03102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07225__A1 (.I(_03102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07207__A1 (.I(_03102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07153__A1 (.I(_03102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07135__A1 (.I(_03102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07117__A1 (.I(_03102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07099__A1 (.I(_03102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07081__A1 (.I(_03102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07063__A1 (.I(_03102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07045__A1 (.I(_03102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07009__A1 (.I(_03102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06991__A1 (.I(_03102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06973__A1 (.I(_03102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06955__A1 (.I(_03102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06937__A1 (.I(_03102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06913__A1 (.I(_03102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07245__A1 (.I(_03104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07227__A1 (.I(_03104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07209__A1 (.I(_03104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07155__A1 (.I(_03104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07137__A1 (.I(_03104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07119__A1 (.I(_03104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07101__A1 (.I(_03104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07083__A1 (.I(_03104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07065__A1 (.I(_03104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07047__A1 (.I(_03104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07011__A1 (.I(_03104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06993__A1 (.I(_03104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06975__A1 (.I(_03104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06957__A1 (.I(_03104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06939__A1 (.I(_03104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06916__A1 (.I(_03104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07247__A1 (.I(_03106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07229__A1 (.I(_03106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07211__A1 (.I(_03106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07157__A1 (.I(_03106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07139__A1 (.I(_03106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07121__A1 (.I(_03106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07103__A1 (.I(_03106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07085__A1 (.I(_03106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07067__A1 (.I(_03106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07049__A1 (.I(_03106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07013__A1 (.I(_03106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06995__A1 (.I(_03106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06977__A1 (.I(_03106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06959__A1 (.I(_03106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06941__A1 (.I(_03106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06919__A1 (.I(_03106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07249__A1 (.I(_03108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07231__A1 (.I(_03108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07213__A1 (.I(_03108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07159__A1 (.I(_03108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07141__A1 (.I(_03108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07123__A1 (.I(_03108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07105__A1 (.I(_03108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07087__A1 (.I(_03108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07069__A1 (.I(_03108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07051__A1 (.I(_03108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07015__A1 (.I(_03108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06997__A1 (.I(_03108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06979__A1 (.I(_03108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06961__A1 (.I(_03108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06943__A1 (.I(_03108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06922__A1 (.I(_03108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07251__A1 (.I(_03110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07233__A1 (.I(_03110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07215__A1 (.I(_03110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07161__A1 (.I(_03110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07143__A1 (.I(_03110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07125__A1 (.I(_03110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07107__A1 (.I(_03110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07089__A1 (.I(_03110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07071__A1 (.I(_03110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07053__A1 (.I(_03110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07017__A1 (.I(_03110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06999__A1 (.I(_03110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06981__A1 (.I(_03110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06963__A1 (.I(_03110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06945__A1 (.I(_03110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06925__A1 (.I(_03110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07253__A1 (.I(_03112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07235__A1 (.I(_03112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07217__A1 (.I(_03112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07163__A1 (.I(_03112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07145__A1 (.I(_03112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07127__A1 (.I(_03112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07109__A1 (.I(_03112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07091__A1 (.I(_03112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07073__A1 (.I(_03112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07055__A1 (.I(_03112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07019__A1 (.I(_03112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07001__A1 (.I(_03112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06983__A1 (.I(_03112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06965__A1 (.I(_03112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06947__A1 (.I(_03112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06928__A1 (.I(_03112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07255__A1 (.I(_03114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07237__A1 (.I(_03114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07219__A1 (.I(_03114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07165__A1 (.I(_03114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07147__A1 (.I(_03114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07129__A1 (.I(_03114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07111__A1 (.I(_03114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07093__A1 (.I(_03114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07075__A1 (.I(_03114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07057__A1 (.I(_03114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07021__A1 (.I(_03114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07003__A1 (.I(_03114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06985__A1 (.I(_03114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06967__A1 (.I(_03114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06949__A1 (.I(_03114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06931__A1 (.I(_03114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06949__A2 (.I(_03117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06948__A2 (.I(_03117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06947__A2 (.I(_03117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06946__A2 (.I(_03117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06945__A2 (.I(_03117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06944__A2 (.I(_03117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06943__A2 (.I(_03117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06942__A2 (.I(_03117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06941__A2 (.I(_03117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06940__A2 (.I(_03117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06939__A2 (.I(_03117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06938__A2 (.I(_03117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06937__A2 (.I(_03117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06936__A2 (.I(_03117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06935__A2 (.I(_03117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06934__A2 (.I(_03117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06967__A2 (.I(_03127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06966__A2 (.I(_03127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06965__A2 (.I(_03127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06964__A2 (.I(_03127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06963__A2 (.I(_03127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06962__A2 (.I(_03127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06961__A2 (.I(_03127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06960__A2 (.I(_03127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06959__A2 (.I(_03127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06958__A2 (.I(_03127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06957__A2 (.I(_03127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06956__A2 (.I(_03127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06955__A2 (.I(_03127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06954__A2 (.I(_03127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06953__A2 (.I(_03127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06952__A2 (.I(_03127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06985__A2 (.I(_03137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06984__A2 (.I(_03137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06983__A2 (.I(_03137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06982__A2 (.I(_03137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06981__A2 (.I(_03137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06980__A2 (.I(_03137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06979__A2 (.I(_03137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06978__A2 (.I(_03137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06977__A2 (.I(_03137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06976__A2 (.I(_03137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06975__A2 (.I(_03137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06974__A2 (.I(_03137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06973__A2 (.I(_03137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06972__A2 (.I(_03137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06971__A2 (.I(_03137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06970__A2 (.I(_03137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07003__A2 (.I(_03147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07002__A2 (.I(_03147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07001__A2 (.I(_03147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07000__A2 (.I(_03147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06999__A2 (.I(_03147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06998__A2 (.I(_03147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06997__A2 (.I(_03147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06996__A2 (.I(_03147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06995__A2 (.I(_03147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06994__A2 (.I(_03147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06993__A2 (.I(_03147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06992__A2 (.I(_03147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06991__A2 (.I(_03147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06990__A2 (.I(_03147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06989__A2 (.I(_03147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06988__A2 (.I(_03147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07021__A2 (.I(_03157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07020__A2 (.I(_03157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07019__A2 (.I(_03157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07018__A2 (.I(_03157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07017__A2 (.I(_03157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07016__A2 (.I(_03157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07015__A2 (.I(_03157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07014__A2 (.I(_03157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07013__A2 (.I(_03157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07012__A2 (.I(_03157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07011__A2 (.I(_03157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07010__A2 (.I(_03157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07009__A2 (.I(_03157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07008__A2 (.I(_03157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07007__A2 (.I(_03157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07006__A2 (.I(_03157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07039__A2 (.I(_03167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07038__A2 (.I(_03167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07037__A2 (.I(_03167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07036__A2 (.I(_03167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07035__A2 (.I(_03167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07034__A2 (.I(_03167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07033__A2 (.I(_03167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07032__A2 (.I(_03167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07031__A2 (.I(_03167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07030__A2 (.I(_03167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07029__A2 (.I(_03167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07028__A2 (.I(_03167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07027__A2 (.I(_03167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07026__A2 (.I(_03167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07025__A2 (.I(_03167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07024__A2 (.I(_03167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07057__A2 (.I(_03177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07056__A2 (.I(_03177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07055__A2 (.I(_03177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07054__A2 (.I(_03177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07053__A2 (.I(_03177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07052__A2 (.I(_03177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07051__A2 (.I(_03177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07050__A2 (.I(_03177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07049__A2 (.I(_03177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07048__A2 (.I(_03177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07047__A2 (.I(_03177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07046__A2 (.I(_03177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07045__A2 (.I(_03177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07044__A2 (.I(_03177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07043__A2 (.I(_03177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07042__A2 (.I(_03177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07075__A2 (.I(_03187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07074__A2 (.I(_03187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07073__A2 (.I(_03187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07072__A2 (.I(_03187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07071__A2 (.I(_03187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07070__A2 (.I(_03187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07069__A2 (.I(_03187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07068__A2 (.I(_03187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07067__A2 (.I(_03187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07066__A2 (.I(_03187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07065__A2 (.I(_03187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07064__A2 (.I(_03187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07063__A2 (.I(_03187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07062__A2 (.I(_03187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07061__A2 (.I(_03187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07060__A2 (.I(_03187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07093__A2 (.I(_03197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07092__A2 (.I(_03197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07091__A2 (.I(_03197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07090__A2 (.I(_03197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07089__A2 (.I(_03197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07088__A2 (.I(_03197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07087__A2 (.I(_03197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07086__A2 (.I(_03197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07085__A2 (.I(_03197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07084__A2 (.I(_03197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07083__A2 (.I(_03197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07082__A2 (.I(_03197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07081__A2 (.I(_03197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07080__A2 (.I(_03197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07079__A2 (.I(_03197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07078__A2 (.I(_03197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07111__A2 (.I(_03207_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07110__A2 (.I(_03207_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07109__A2 (.I(_03207_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07108__A2 (.I(_03207_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07107__A2 (.I(_03207_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07106__A2 (.I(_03207_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07105__A2 (.I(_03207_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07104__A2 (.I(_03207_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07103__A2 (.I(_03207_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07102__A2 (.I(_03207_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07101__A2 (.I(_03207_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07100__A2 (.I(_03207_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07099__A2 (.I(_03207_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07098__A2 (.I(_03207_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07097__A2 (.I(_03207_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07096__A2 (.I(_03207_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07129__A2 (.I(_03217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07128__A2 (.I(_03217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07127__A2 (.I(_03217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07126__A2 (.I(_03217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07125__A2 (.I(_03217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07124__A2 (.I(_03217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07123__A2 (.I(_03217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07122__A2 (.I(_03217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07121__A2 (.I(_03217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07120__A2 (.I(_03217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07119__A2 (.I(_03217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07118__A2 (.I(_03217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07117__A2 (.I(_03217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07116__A2 (.I(_03217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07115__A2 (.I(_03217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07114__A2 (.I(_03217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07147__A2 (.I(_03227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07146__A2 (.I(_03227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07145__A2 (.I(_03227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07144__A2 (.I(_03227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07143__A2 (.I(_03227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07142__A2 (.I(_03227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07141__A2 (.I(_03227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07140__A2 (.I(_03227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07139__A2 (.I(_03227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07138__A2 (.I(_03227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07137__A2 (.I(_03227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07136__A2 (.I(_03227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07135__A2 (.I(_03227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07134__A2 (.I(_03227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07133__A2 (.I(_03227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07132__A2 (.I(_03227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07165__A2 (.I(_03237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07164__A2 (.I(_03237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07163__A2 (.I(_03237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07162__A2 (.I(_03237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07161__A2 (.I(_03237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07160__A2 (.I(_03237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07159__A2 (.I(_03237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07158__A2 (.I(_03237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07157__A2 (.I(_03237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07156__A2 (.I(_03237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07155__A2 (.I(_03237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07154__A2 (.I(_03237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07153__A2 (.I(_03237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07152__A2 (.I(_03237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07151__A2 (.I(_03237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07150__A2 (.I(_03237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07183__A2 (.I(_03247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07182__A2 (.I(_03247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07181__A2 (.I(_03247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07180__A2 (.I(_03247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07179__A2 (.I(_03247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07178__A2 (.I(_03247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07177__A2 (.I(_03247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07176__A2 (.I(_03247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07175__A2 (.I(_03247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07174__A2 (.I(_03247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07173__A2 (.I(_03247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07172__A2 (.I(_03247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07171__A2 (.I(_03247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07170__A2 (.I(_03247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07169__A2 (.I(_03247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07168__A2 (.I(_03247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07201__A2 (.I(_03257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07200__A2 (.I(_03257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07199__A2 (.I(_03257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07198__A2 (.I(_03257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07197__A2 (.I(_03257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07196__A2 (.I(_03257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07195__A2 (.I(_03257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07194__A2 (.I(_03257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07193__A2 (.I(_03257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07192__A2 (.I(_03257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07191__A2 (.I(_03257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07190__A2 (.I(_03257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07189__A2 (.I(_03257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07188__A2 (.I(_03257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07187__A2 (.I(_03257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07186__A2 (.I(_03257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07219__A2 (.I(_03267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07218__A2 (.I(_03267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07217__A2 (.I(_03267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07216__A2 (.I(_03267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07215__A2 (.I(_03267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07214__A2 (.I(_03267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07213__A2 (.I(_03267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07212__A2 (.I(_03267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07211__A2 (.I(_03267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07210__A2 (.I(_03267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07209__A2 (.I(_03267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07208__A2 (.I(_03267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07207__A2 (.I(_03267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07206__A2 (.I(_03267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07205__A2 (.I(_03267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07204__A2 (.I(_03267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07237__A2 (.I(_03277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07236__A2 (.I(_03277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07235__A2 (.I(_03277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07234__A2 (.I(_03277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07233__A2 (.I(_03277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07232__A2 (.I(_03277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07231__A2 (.I(_03277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07230__A2 (.I(_03277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07229__A2 (.I(_03277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07228__A2 (.I(_03277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07227__A2 (.I(_03277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07226__A2 (.I(_03277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07225__A2 (.I(_03277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07224__A2 (.I(_03277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07223__A2 (.I(_03277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07222__A2 (.I(_03277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07255__A2 (.I(_03287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07254__A2 (.I(_03287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07253__A2 (.I(_03287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07252__A2 (.I(_03287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07251__A2 (.I(_03287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07250__A2 (.I(_03287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07249__A2 (.I(_03287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07248__A2 (.I(_03287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07247__A2 (.I(_03287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07246__A2 (.I(_03287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07245__A2 (.I(_03287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07244__A2 (.I(_03287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07243__A2 (.I(_03287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07242__A2 (.I(_03287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07241__A2 (.I(_03287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07240__A2 (.I(_03287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07273__A2 (.I(_03297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07272__A2 (.I(_03297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07271__A2 (.I(_03297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07270__A2 (.I(_03297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07269__A2 (.I(_03297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07268__A2 (.I(_03297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07267__A2 (.I(_03297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07266__A2 (.I(_03297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07265__A2 (.I(_03297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07264__A2 (.I(_03297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07263__A2 (.I(_03297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07262__A2 (.I(_03297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07261__A2 (.I(_03297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07260__A2 (.I(_03297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07259__A2 (.I(_03297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07258__A2 (.I(_03297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07573__A1 (.I(_03306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07555__A1 (.I(_03306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07537__A1 (.I(_03306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07519__A1 (.I(_03306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07501__A1 (.I(_03306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07483__A1 (.I(_03306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07465__A1 (.I(_03306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07447__A1 (.I(_03306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07429__A1 (.I(_03306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07411__A1 (.I(_03306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07393__A1 (.I(_03306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07357__A1 (.I(_03306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07339__A1 (.I(_03306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07321__A1 (.I(_03306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07303__A1 (.I(_03306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07278__A1 (.I(_03306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07299__A2 (.I(_03308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07298__A2 (.I(_03308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07296__A2 (.I(_03308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07295__A2 (.I(_03308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07293__A2 (.I(_03308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07292__A2 (.I(_03308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07290__A2 (.I(_03308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07289__A2 (.I(_03308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07287__A2 (.I(_03308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07286__A2 (.I(_03308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07284__A2 (.I(_03308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07283__A2 (.I(_03308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07281__A2 (.I(_03308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07280__A2 (.I(_03308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07278__A2 (.I(_03308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07277__A2 (.I(_03308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07575__A1 (.I(_03310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07557__A1 (.I(_03310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07539__A1 (.I(_03310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07521__A1 (.I(_03310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07503__A1 (.I(_03310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07485__A1 (.I(_03310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07467__A1 (.I(_03310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07449__A1 (.I(_03310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07431__A1 (.I(_03310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07413__A1 (.I(_03310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07395__A1 (.I(_03310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07359__A1 (.I(_03310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07341__A1 (.I(_03310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07323__A1 (.I(_03310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07305__A1 (.I(_03310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07281__A1 (.I(_03310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07577__A1 (.I(_03312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07559__A1 (.I(_03312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07541__A1 (.I(_03312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07523__A1 (.I(_03312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07505__A1 (.I(_03312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07487__A1 (.I(_03312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07469__A1 (.I(_03312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07451__A1 (.I(_03312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07433__A1 (.I(_03312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07415__A1 (.I(_03312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07397__A1 (.I(_03312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07361__A1 (.I(_03312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07343__A1 (.I(_03312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07325__A1 (.I(_03312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07307__A1 (.I(_03312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07284__A1 (.I(_03312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07579__A1 (.I(_03314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07561__A1 (.I(_03314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07543__A1 (.I(_03314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07525__A1 (.I(_03314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07507__A1 (.I(_03314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07489__A1 (.I(_03314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07471__A1 (.I(_03314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07453__A1 (.I(_03314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07435__A1 (.I(_03314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07417__A1 (.I(_03314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07399__A1 (.I(_03314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07363__A1 (.I(_03314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07345__A1 (.I(_03314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07327__A1 (.I(_03314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07309__A1 (.I(_03314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07287__A1 (.I(_03314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07581__A1 (.I(_03316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07563__A1 (.I(_03316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07545__A1 (.I(_03316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07527__A1 (.I(_03316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07509__A1 (.I(_03316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07491__A1 (.I(_03316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07473__A1 (.I(_03316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07455__A1 (.I(_03316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07437__A1 (.I(_03316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07419__A1 (.I(_03316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07401__A1 (.I(_03316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07365__A1 (.I(_03316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07347__A1 (.I(_03316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07329__A1 (.I(_03316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07311__A1 (.I(_03316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07290__A1 (.I(_03316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07583__A1 (.I(_03318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07565__A1 (.I(_03318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07547__A1 (.I(_03318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07529__A1 (.I(_03318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07511__A1 (.I(_03318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07493__A1 (.I(_03318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07475__A1 (.I(_03318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07457__A1 (.I(_03318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07439__A1 (.I(_03318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07421__A1 (.I(_03318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07403__A1 (.I(_03318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07367__A1 (.I(_03318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07349__A1 (.I(_03318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07331__A1 (.I(_03318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07313__A1 (.I(_03318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07293__A1 (.I(_03318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07585__A1 (.I(_03320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07567__A1 (.I(_03320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07549__A1 (.I(_03320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07531__A1 (.I(_03320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07513__A1 (.I(_03320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07495__A1 (.I(_03320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07477__A1 (.I(_03320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07459__A1 (.I(_03320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07441__A1 (.I(_03320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07423__A1 (.I(_03320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07405__A1 (.I(_03320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07369__A1 (.I(_03320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07351__A1 (.I(_03320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07333__A1 (.I(_03320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07315__A1 (.I(_03320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07296__A1 (.I(_03320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07587__A1 (.I(_03322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07569__A1 (.I(_03322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07551__A1 (.I(_03322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07533__A1 (.I(_03322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07515__A1 (.I(_03322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07497__A1 (.I(_03322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07479__A1 (.I(_03322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07461__A1 (.I(_03322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07443__A1 (.I(_03322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07425__A1 (.I(_03322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07407__A1 (.I(_03322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07371__A1 (.I(_03322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07353__A1 (.I(_03322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07335__A1 (.I(_03322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07317__A1 (.I(_03322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07299__A1 (.I(_03322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07317__A2 (.I(_03325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07316__A2 (.I(_03325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07315__A2 (.I(_03325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07314__A2 (.I(_03325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07313__A2 (.I(_03325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07312__A2 (.I(_03325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07311__A2 (.I(_03325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07310__A2 (.I(_03325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07309__A2 (.I(_03325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07308__A2 (.I(_03325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07307__A2 (.I(_03325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07306__A2 (.I(_03325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07305__A2 (.I(_03325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07304__A2 (.I(_03325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07303__A2 (.I(_03325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07302__A2 (.I(_03325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07335__A2 (.I(_03335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07334__A2 (.I(_03335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07333__A2 (.I(_03335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07332__A2 (.I(_03335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07331__A2 (.I(_03335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07330__A2 (.I(_03335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07329__A2 (.I(_03335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07328__A2 (.I(_03335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07327__A2 (.I(_03335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07326__A2 (.I(_03335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07325__A2 (.I(_03335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07324__A2 (.I(_03335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07323__A2 (.I(_03335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07322__A2 (.I(_03335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07321__A2 (.I(_03335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07320__A2 (.I(_03335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07353__A2 (.I(_03345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07352__A2 (.I(_03345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07351__A2 (.I(_03345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07350__A2 (.I(_03345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07349__A2 (.I(_03345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07348__A2 (.I(_03345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07347__A2 (.I(_03345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07346__A2 (.I(_03345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07345__A2 (.I(_03345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07344__A2 (.I(_03345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07343__A2 (.I(_03345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07342__A2 (.I(_03345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07341__A2 (.I(_03345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07340__A2 (.I(_03345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07339__A2 (.I(_03345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07338__A2 (.I(_03345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07371__A2 (.I(_03355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07370__A2 (.I(_03355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07369__A2 (.I(_03355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07368__A2 (.I(_03355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07367__A2 (.I(_03355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07366__A2 (.I(_03355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07365__A2 (.I(_03355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07364__A2 (.I(_03355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07363__A2 (.I(_03355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07362__A2 (.I(_03355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07361__A2 (.I(_03355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07360__A2 (.I(_03355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07359__A2 (.I(_03355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07358__A2 (.I(_03355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07357__A2 (.I(_03355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07356__A2 (.I(_03355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07389__A2 (.I(_03365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07388__A2 (.I(_03365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07387__A2 (.I(_03365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07386__A2 (.I(_03365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07385__A2 (.I(_03365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07384__A2 (.I(_03365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07383__A2 (.I(_03365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07382__A2 (.I(_03365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07381__A2 (.I(_03365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07380__A2 (.I(_03365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07379__A2 (.I(_03365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07378__A2 (.I(_03365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07377__A2 (.I(_03365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07376__A2 (.I(_03365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07375__A2 (.I(_03365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07374__A2 (.I(_03365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07407__A2 (.I(_03375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07406__A2 (.I(_03375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07405__A2 (.I(_03375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07404__A2 (.I(_03375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07403__A2 (.I(_03375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07402__A2 (.I(_03375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07401__A2 (.I(_03375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07400__A2 (.I(_03375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07399__A2 (.I(_03375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07398__A2 (.I(_03375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07397__A2 (.I(_03375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07396__A2 (.I(_03375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07395__A2 (.I(_03375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07394__A2 (.I(_03375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07393__A2 (.I(_03375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07392__A2 (.I(_03375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07425__A2 (.I(_03385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07424__A2 (.I(_03385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07423__A2 (.I(_03385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07422__A2 (.I(_03385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07421__A2 (.I(_03385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07420__A2 (.I(_03385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07419__A2 (.I(_03385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07418__A2 (.I(_03385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07417__A2 (.I(_03385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07416__A2 (.I(_03385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07415__A2 (.I(_03385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07414__A2 (.I(_03385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07413__A2 (.I(_03385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07412__A2 (.I(_03385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07411__A2 (.I(_03385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07410__A2 (.I(_03385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07443__A2 (.I(_03395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07442__A2 (.I(_03395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07441__A2 (.I(_03395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07440__A2 (.I(_03395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07439__A2 (.I(_03395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07438__A2 (.I(_03395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07437__A2 (.I(_03395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07436__A2 (.I(_03395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07435__A2 (.I(_03395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07434__A2 (.I(_03395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07433__A2 (.I(_03395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07432__A2 (.I(_03395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07431__A2 (.I(_03395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07430__A2 (.I(_03395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07429__A2 (.I(_03395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07428__A2 (.I(_03395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07461__A2 (.I(_03405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07460__A2 (.I(_03405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07459__A2 (.I(_03405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07458__A2 (.I(_03405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07457__A2 (.I(_03405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07456__A2 (.I(_03405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07455__A2 (.I(_03405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07454__A2 (.I(_03405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07453__A2 (.I(_03405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07452__A2 (.I(_03405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07451__A2 (.I(_03405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07450__A2 (.I(_03405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07449__A2 (.I(_03405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07448__A2 (.I(_03405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07447__A2 (.I(_03405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07446__A2 (.I(_03405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07479__A2 (.I(_03415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07478__A2 (.I(_03415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07477__A2 (.I(_03415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07476__A2 (.I(_03415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07475__A2 (.I(_03415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07474__A2 (.I(_03415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07473__A2 (.I(_03415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07472__A2 (.I(_03415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07471__A2 (.I(_03415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07470__A2 (.I(_03415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07469__A2 (.I(_03415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07468__A2 (.I(_03415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07467__A2 (.I(_03415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07466__A2 (.I(_03415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07465__A2 (.I(_03415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07464__A2 (.I(_03415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07497__A2 (.I(_03425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07496__A2 (.I(_03425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07495__A2 (.I(_03425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07494__A2 (.I(_03425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07493__A2 (.I(_03425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07492__A2 (.I(_03425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07491__A2 (.I(_03425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07490__A2 (.I(_03425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07489__A2 (.I(_03425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07488__A2 (.I(_03425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07487__A2 (.I(_03425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07486__A2 (.I(_03425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07485__A2 (.I(_03425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07484__A2 (.I(_03425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07483__A2 (.I(_03425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07482__A2 (.I(_03425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07515__A2 (.I(_03435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07514__A2 (.I(_03435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07513__A2 (.I(_03435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07512__A2 (.I(_03435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07511__A2 (.I(_03435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07510__A2 (.I(_03435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07509__A2 (.I(_03435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07508__A2 (.I(_03435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07507__A2 (.I(_03435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07506__A2 (.I(_03435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07505__A2 (.I(_03435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07504__A2 (.I(_03435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07503__A2 (.I(_03435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07502__A2 (.I(_03435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07501__A2 (.I(_03435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07500__A2 (.I(_03435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07533__A2 (.I(_03445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07532__A2 (.I(_03445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07531__A2 (.I(_03445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07530__A2 (.I(_03445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07529__A2 (.I(_03445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07528__A2 (.I(_03445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07527__A2 (.I(_03445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07526__A2 (.I(_03445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07525__A2 (.I(_03445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07524__A2 (.I(_03445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07523__A2 (.I(_03445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07522__A2 (.I(_03445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07521__A2 (.I(_03445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07520__A2 (.I(_03445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07519__A2 (.I(_03445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07518__A2 (.I(_03445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07551__A2 (.I(_03455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07550__A2 (.I(_03455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07549__A2 (.I(_03455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07548__A2 (.I(_03455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07547__A2 (.I(_03455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07546__A2 (.I(_03455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07545__A2 (.I(_03455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07544__A2 (.I(_03455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07543__A2 (.I(_03455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07542__A2 (.I(_03455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07541__A2 (.I(_03455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07540__A2 (.I(_03455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07539__A2 (.I(_03455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07538__A2 (.I(_03455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07537__A2 (.I(_03455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07536__A2 (.I(_03455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07569__A2 (.I(_03465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07568__A2 (.I(_03465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07567__A2 (.I(_03465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07566__A2 (.I(_03465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07565__A2 (.I(_03465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07564__A2 (.I(_03465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07563__A2 (.I(_03465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07562__A2 (.I(_03465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07561__A2 (.I(_03465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07560__A2 (.I(_03465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07559__A2 (.I(_03465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07558__A2 (.I(_03465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07557__A2 (.I(_03465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07556__A2 (.I(_03465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07555__A2 (.I(_03465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07554__A2 (.I(_03465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07587__A2 (.I(_03475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07586__A2 (.I(_03475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07585__A2 (.I(_03475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07584__A2 (.I(_03475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07583__A2 (.I(_03475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07582__A2 (.I(_03475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07581__A2 (.I(_03475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07580__A2 (.I(_03475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07579__A2 (.I(_03475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07578__A2 (.I(_03475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07577__A2 (.I(_03475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07576__A2 (.I(_03475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07575__A2 (.I(_03475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07574__A2 (.I(_03475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07573__A2 (.I(_03475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07572__A2 (.I(_03475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07605__A2 (.I(_03485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07604__A2 (.I(_03485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07603__A2 (.I(_03485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07602__A2 (.I(_03485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07601__A2 (.I(_03485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07600__A2 (.I(_03485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07599__A2 (.I(_03485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07598__A2 (.I(_03485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07597__A2 (.I(_03485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07596__A2 (.I(_03485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07595__A2 (.I(_03485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07594__A2 (.I(_03485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07593__A2 (.I(_03485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07592__A2 (.I(_03485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07591__A2 (.I(_03485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07590__A2 (.I(_03485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07928__A1 (.I(_03494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07910__A1 (.I(_03494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07892__A1 (.I(_03494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07874__A1 (.I(_03494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07836__A1 (.I(_03494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07818__A1 (.I(_03494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07779__A1 (.I(_03494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07761__A1 (.I(_03494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07743__A1 (.I(_03494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07725__A1 (.I(_03494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07707__A1 (.I(_03494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07689__A1 (.I(_03494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07671__A1 (.I(_03494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07653__A1 (.I(_03494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07635__A1 (.I(_03494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07610__A1 (.I(_03494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07631__A2 (.I(_03496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07630__A2 (.I(_03496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07628__A2 (.I(_03496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07627__A2 (.I(_03496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07625__A2 (.I(_03496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07624__A2 (.I(_03496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07622__A2 (.I(_03496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07621__A2 (.I(_03496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07619__A2 (.I(_03496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07618__A2 (.I(_03496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07616__A2 (.I(_03496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07615__A2 (.I(_03496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07613__A2 (.I(_03496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07612__A2 (.I(_03496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07610__A2 (.I(_03496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07609__A2 (.I(_03496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07930__A1 (.I(_03498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07912__A1 (.I(_03498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07894__A1 (.I(_03498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07876__A1 (.I(_03498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07838__A1 (.I(_03498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07820__A1 (.I(_03498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07781__A1 (.I(_03498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07763__A1 (.I(_03498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07745__A1 (.I(_03498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07727__A1 (.I(_03498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07709__A1 (.I(_03498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07691__A1 (.I(_03498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07673__A1 (.I(_03498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07655__A1 (.I(_03498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07637__A1 (.I(_03498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07613__A1 (.I(_03498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07932__A1 (.I(_03500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07914__A1 (.I(_03500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07896__A1 (.I(_03500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07878__A1 (.I(_03500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07840__A1 (.I(_03500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07822__A1 (.I(_03500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07783__A1 (.I(_03500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07765__A1 (.I(_03500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07747__A1 (.I(_03500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07729__A1 (.I(_03500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07711__A1 (.I(_03500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07693__A1 (.I(_03500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07675__A1 (.I(_03500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07657__A1 (.I(_03500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07639__A1 (.I(_03500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07616__A1 (.I(_03500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07934__A1 (.I(_03502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07916__A1 (.I(_03502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07898__A1 (.I(_03502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07880__A1 (.I(_03502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07842__A1 (.I(_03502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07824__A1 (.I(_03502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07785__A1 (.I(_03502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07767__A1 (.I(_03502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07749__A1 (.I(_03502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07731__A1 (.I(_03502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07713__A1 (.I(_03502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07695__A1 (.I(_03502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07677__A1 (.I(_03502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07659__A1 (.I(_03502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07641__A1 (.I(_03502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07619__A1 (.I(_03502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07936__A1 (.I(_03504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07918__A1 (.I(_03504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07900__A1 (.I(_03504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07882__A1 (.I(_03504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07844__A1 (.I(_03504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07826__A1 (.I(_03504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07787__A1 (.I(_03504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07769__A1 (.I(_03504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07751__A1 (.I(_03504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07733__A1 (.I(_03504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07715__A1 (.I(_03504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07697__A1 (.I(_03504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07679__A1 (.I(_03504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07661__A1 (.I(_03504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07643__A1 (.I(_03504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07622__A1 (.I(_03504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07938__A1 (.I(_03506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07920__A1 (.I(_03506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07902__A1 (.I(_03506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07884__A1 (.I(_03506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07846__A1 (.I(_03506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07828__A1 (.I(_03506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07789__A1 (.I(_03506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07771__A1 (.I(_03506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07753__A1 (.I(_03506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07735__A1 (.I(_03506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07717__A1 (.I(_03506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07699__A1 (.I(_03506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07681__A1 (.I(_03506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07663__A1 (.I(_03506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07645__A1 (.I(_03506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07625__A1 (.I(_03506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07940__A1 (.I(_03508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07922__A1 (.I(_03508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07904__A1 (.I(_03508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07886__A1 (.I(_03508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07848__A1 (.I(_03508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07830__A1 (.I(_03508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07791__A1 (.I(_03508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07773__A1 (.I(_03508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07755__A1 (.I(_03508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07737__A1 (.I(_03508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07719__A1 (.I(_03508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07701__A1 (.I(_03508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07683__A1 (.I(_03508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07665__A1 (.I(_03508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07647__A1 (.I(_03508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07628__A1 (.I(_03508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07942__A1 (.I(_03510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07924__A1 (.I(_03510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07906__A1 (.I(_03510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07888__A1 (.I(_03510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07850__A1 (.I(_03510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07832__A1 (.I(_03510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07793__A1 (.I(_03510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07775__A1 (.I(_03510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07757__A1 (.I(_03510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07739__A1 (.I(_03510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07721__A1 (.I(_03510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07703__A1 (.I(_03510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07685__A1 (.I(_03510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07667__A1 (.I(_03510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07649__A1 (.I(_03510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07631__A1 (.I(_03510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07649__A2 (.I(_03513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07648__A2 (.I(_03513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07647__A2 (.I(_03513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07646__A2 (.I(_03513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07645__A2 (.I(_03513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07644__A2 (.I(_03513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07643__A2 (.I(_03513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07642__A2 (.I(_03513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07641__A2 (.I(_03513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07640__A2 (.I(_03513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07639__A2 (.I(_03513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07638__A2 (.I(_03513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07637__A2 (.I(_03513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07636__A2 (.I(_03513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07635__A2 (.I(_03513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07634__A2 (.I(_03513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07667__A2 (.I(_03523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07666__A2 (.I(_03523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07665__A2 (.I(_03523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07664__A2 (.I(_03523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07663__A2 (.I(_03523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07662__A2 (.I(_03523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07661__A2 (.I(_03523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07660__A2 (.I(_03523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07659__A2 (.I(_03523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07658__A2 (.I(_03523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07657__A2 (.I(_03523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07656__A2 (.I(_03523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07655__A2 (.I(_03523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07654__A2 (.I(_03523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07653__A2 (.I(_03523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07652__A2 (.I(_03523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07685__A2 (.I(_03533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07684__A2 (.I(_03533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07683__A2 (.I(_03533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07682__A2 (.I(_03533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07681__A2 (.I(_03533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07680__A2 (.I(_03533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07679__A2 (.I(_03533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07678__A2 (.I(_03533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07677__A2 (.I(_03533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07676__A2 (.I(_03533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07675__A2 (.I(_03533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07674__A2 (.I(_03533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07673__A2 (.I(_03533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07672__A2 (.I(_03533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07671__A2 (.I(_03533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07670__A2 (.I(_03533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07703__A2 (.I(_03543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07702__A2 (.I(_03543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07701__A2 (.I(_03543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07700__A2 (.I(_03543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07699__A2 (.I(_03543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07698__A2 (.I(_03543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07697__A2 (.I(_03543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07696__A2 (.I(_03543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07695__A2 (.I(_03543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07694__A2 (.I(_03543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07693__A2 (.I(_03543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07692__A2 (.I(_03543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07691__A2 (.I(_03543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07690__A2 (.I(_03543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07689__A2 (.I(_03543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07688__A2 (.I(_03543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07721__A2 (.I(_03553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07720__A2 (.I(_03553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07719__A2 (.I(_03553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07718__A2 (.I(_03553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07717__A2 (.I(_03553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07716__A2 (.I(_03553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07715__A2 (.I(_03553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07714__A2 (.I(_03553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07713__A2 (.I(_03553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07712__A2 (.I(_03553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07711__A2 (.I(_03553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07710__A2 (.I(_03553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07709__A2 (.I(_03553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07708__A2 (.I(_03553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07707__A2 (.I(_03553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07706__A2 (.I(_03553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07739__A2 (.I(_03563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07738__A2 (.I(_03563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07737__A2 (.I(_03563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07736__A2 (.I(_03563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07735__A2 (.I(_03563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07734__A2 (.I(_03563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07733__A2 (.I(_03563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07732__A2 (.I(_03563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07731__A2 (.I(_03563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07730__A2 (.I(_03563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07729__A2 (.I(_03563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07728__A2 (.I(_03563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07727__A2 (.I(_03563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07726__A2 (.I(_03563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07725__A2 (.I(_03563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07724__A2 (.I(_03563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07757__A2 (.I(_03573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07756__A2 (.I(_03573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07755__A2 (.I(_03573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07754__A2 (.I(_03573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07753__A2 (.I(_03573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07752__A2 (.I(_03573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07751__A2 (.I(_03573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07750__A2 (.I(_03573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07749__A2 (.I(_03573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07748__A2 (.I(_03573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07747__A2 (.I(_03573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07746__A2 (.I(_03573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07745__A2 (.I(_03573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07744__A2 (.I(_03573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07743__A2 (.I(_03573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07742__A2 (.I(_03573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07775__A2 (.I(_03583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07774__A2 (.I(_03583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07773__A2 (.I(_03583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07772__A2 (.I(_03583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07771__A2 (.I(_03583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07770__A2 (.I(_03583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07769__A2 (.I(_03583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07768__A2 (.I(_03583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07767__A2 (.I(_03583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07766__A2 (.I(_03583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07765__A2 (.I(_03583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07764__A2 (.I(_03583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07763__A2 (.I(_03583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07762__A2 (.I(_03583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07761__A2 (.I(_03583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07760__A2 (.I(_03583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07793__A2 (.I(_03593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07792__A2 (.I(_03593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07791__A2 (.I(_03593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07790__A2 (.I(_03593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07789__A2 (.I(_03593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07788__A2 (.I(_03593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07787__A2 (.I(_03593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07786__A2 (.I(_03593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07785__A2 (.I(_03593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07784__A2 (.I(_03593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07783__A2 (.I(_03593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07782__A2 (.I(_03593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07781__A2 (.I(_03593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07780__A2 (.I(_03593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07779__A2 (.I(_03593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07778__A2 (.I(_03593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09516__A2 (.I(_03605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07802__A2 (.I(_03605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07801__A2 (.I(_03605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07800__A2 (.I(_03605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07799__A3 (.I(_03605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09690__A2 (.I(_03611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09526__A2 (.I(_03611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07869__A2 (.I(_03611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07854__A2 (.I(_03611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07852__A2 (.I(_03611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07808__A2 (.I(_03611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07832__A2 (.I(_03616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07831__A2 (.I(_03616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07830__A2 (.I(_03616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07829__A2 (.I(_03616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07828__A2 (.I(_03616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07827__A2 (.I(_03616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07826__A2 (.I(_03616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07825__A2 (.I(_03616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07824__A2 (.I(_03616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07823__A2 (.I(_03616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07822__A2 (.I(_03616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07821__A2 (.I(_03616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07820__A2 (.I(_03616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07819__A2 (.I(_03616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07818__A2 (.I(_03616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07817__A2 (.I(_03616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07850__A2 (.I(_03626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07849__A2 (.I(_03626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07848__A2 (.I(_03626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07847__A2 (.I(_03626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07846__A2 (.I(_03626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07845__A2 (.I(_03626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07844__A2 (.I(_03626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07843__A2 (.I(_03626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07842__A2 (.I(_03626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07841__A2 (.I(_03626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07840__A2 (.I(_03626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07839__A2 (.I(_03626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07838__A2 (.I(_03626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07837__A2 (.I(_03626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07836__A2 (.I(_03626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07835__A2 (.I(_03626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07888__A2 (.I(_03652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07887__A2 (.I(_03652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07886__A2 (.I(_03652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07885__A2 (.I(_03652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07884__A2 (.I(_03652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07883__A2 (.I(_03652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07882__A2 (.I(_03652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07881__A2 (.I(_03652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07880__A2 (.I(_03652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07879__A2 (.I(_03652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07878__A2 (.I(_03652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07877__A2 (.I(_03652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07876__A2 (.I(_03652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07875__A2 (.I(_03652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07874__A2 (.I(_03652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07873__A2 (.I(_03652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07906__A2 (.I(_03662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07905__A2 (.I(_03662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07904__A2 (.I(_03662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07903__A2 (.I(_03662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07902__A2 (.I(_03662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07901__A2 (.I(_03662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07900__A2 (.I(_03662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07899__A2 (.I(_03662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07898__A2 (.I(_03662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07897__A2 (.I(_03662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07896__A2 (.I(_03662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07895__A2 (.I(_03662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07894__A2 (.I(_03662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07893__A2 (.I(_03662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07892__A2 (.I(_03662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07891__A2 (.I(_03662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07924__A2 (.I(_03672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07923__A2 (.I(_03672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07922__A2 (.I(_03672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07921__A2 (.I(_03672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07920__A2 (.I(_03672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07919__A2 (.I(_03672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07918__A2 (.I(_03672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07917__A2 (.I(_03672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07916__A2 (.I(_03672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07915__A2 (.I(_03672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07914__A2 (.I(_03672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07913__A2 (.I(_03672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07912__A2 (.I(_03672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07911__A2 (.I(_03672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07910__A2 (.I(_03672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07909__A2 (.I(_03672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07942__A2 (.I(_03682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07941__A2 (.I(_03682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07940__A2 (.I(_03682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07939__A2 (.I(_03682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07938__A2 (.I(_03682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07937__A2 (.I(_03682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07936__A2 (.I(_03682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07935__A2 (.I(_03682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07934__A2 (.I(_03682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07933__A2 (.I(_03682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07932__A2 (.I(_03682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07931__A2 (.I(_03682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07930__A2 (.I(_03682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07929__A2 (.I(_03682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07928__A2 (.I(_03682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07927__A2 (.I(_03682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08968__A1 (.I(_03691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08911__A1 (.I(_03691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08857__A1 (.I(_03691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08765__A1 (.I(_03691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08672__A1 (.I(_03691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08654__A1 (.I(_03691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08426__A1 (.I(_03691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08251__A1 (.I(_03691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08116__A1 (.I(_03691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08098__A1 (.I(_03691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08080__A1 (.I(_03691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08062__A1 (.I(_03691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08044__A1 (.I(_03691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07990__A1 (.I(_03691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07972__A1 (.I(_03691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07947__A1 (.I(_03691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07968__A2 (.I(_03693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07967__A2 (.I(_03693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07965__A2 (.I(_03693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07964__A2 (.I(_03693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07962__A2 (.I(_03693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07961__A2 (.I(_03693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07959__A2 (.I(_03693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07958__A2 (.I(_03693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07956__A2 (.I(_03693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07955__A2 (.I(_03693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07953__A2 (.I(_03693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07952__A2 (.I(_03693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07950__A2 (.I(_03693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07949__A2 (.I(_03693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07947__A2 (.I(_03693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07946__A2 (.I(_03693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08970__A1 (.I(_03695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08913__A1 (.I(_03695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08859__A1 (.I(_03695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08767__A1 (.I(_03695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08674__A1 (.I(_03695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08656__A1 (.I(_03695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08428__A1 (.I(_03695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08253__A1 (.I(_03695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08118__A1 (.I(_03695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08100__A1 (.I(_03695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08082__A1 (.I(_03695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08064__A1 (.I(_03695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08046__A1 (.I(_03695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07992__A1 (.I(_03695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07974__A1 (.I(_03695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07950__A1 (.I(_03695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08972__A1 (.I(_03697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08915__A1 (.I(_03697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08861__A1 (.I(_03697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08769__A1 (.I(_03697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08676__A1 (.I(_03697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08658__A1 (.I(_03697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08430__A1 (.I(_03697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08255__A1 (.I(_03697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08120__A1 (.I(_03697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08102__A1 (.I(_03697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08084__A1 (.I(_03697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08066__A1 (.I(_03697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08048__A1 (.I(_03697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07994__A1 (.I(_03697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07976__A1 (.I(_03697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07953__A1 (.I(_03697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08974__A1 (.I(_03699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08917__A1 (.I(_03699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08863__A1 (.I(_03699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08771__A1 (.I(_03699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08678__A1 (.I(_03699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08660__A1 (.I(_03699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08432__A1 (.I(_03699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08257__A1 (.I(_03699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08122__A1 (.I(_03699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08104__A1 (.I(_03699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08086__A1 (.I(_03699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08068__A1 (.I(_03699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08050__A1 (.I(_03699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07996__A1 (.I(_03699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07978__A1 (.I(_03699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07956__A1 (.I(_03699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08976__A1 (.I(_03701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08919__A1 (.I(_03701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08865__A1 (.I(_03701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08773__A1 (.I(_03701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08680__A1 (.I(_03701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08662__A1 (.I(_03701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08434__A1 (.I(_03701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08259__A1 (.I(_03701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08124__A1 (.I(_03701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08106__A1 (.I(_03701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08088__A1 (.I(_03701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08070__A1 (.I(_03701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08052__A1 (.I(_03701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07998__A1 (.I(_03701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07980__A1 (.I(_03701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07959__A1 (.I(_03701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08978__A1 (.I(_03703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08921__A1 (.I(_03703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08867__A1 (.I(_03703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08775__A1 (.I(_03703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08682__A1 (.I(_03703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08664__A1 (.I(_03703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08436__A1 (.I(_03703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08261__A1 (.I(_03703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08126__A1 (.I(_03703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08108__A1 (.I(_03703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08090__A1 (.I(_03703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08072__A1 (.I(_03703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08054__A1 (.I(_03703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08000__A1 (.I(_03703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07982__A1 (.I(_03703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07962__A1 (.I(_03703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08980__A1 (.I(_03705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08923__A1 (.I(_03705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08869__A1 (.I(_03705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08777__A1 (.I(_03705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08684__A1 (.I(_03705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08666__A1 (.I(_03705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08438__A1 (.I(_03705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08263__A1 (.I(_03705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08128__A1 (.I(_03705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08110__A1 (.I(_03705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08092__A1 (.I(_03705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08074__A1 (.I(_03705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08056__A1 (.I(_03705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08002__A1 (.I(_03705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07984__A1 (.I(_03705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07965__A1 (.I(_03705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08982__A1 (.I(_03707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08925__A1 (.I(_03707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08871__A1 (.I(_03707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08779__A1 (.I(_03707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08686__A1 (.I(_03707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08668__A1 (.I(_03707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08440__A1 (.I(_03707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08265__A1 (.I(_03707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08130__A1 (.I(_03707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08112__A1 (.I(_03707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08094__A1 (.I(_03707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08076__A1 (.I(_03707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08058__A1 (.I(_03707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08004__A1 (.I(_03707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07986__A1 (.I(_03707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07968__A1 (.I(_03707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07986__A2 (.I(_03710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07985__A2 (.I(_03710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07984__A2 (.I(_03710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07983__A2 (.I(_03710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07982__A2 (.I(_03710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07981__A2 (.I(_03710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07980__A2 (.I(_03710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07979__A2 (.I(_03710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07978__A2 (.I(_03710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07977__A2 (.I(_03710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07976__A2 (.I(_03710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07975__A2 (.I(_03710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07974__A2 (.I(_03710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07973__A2 (.I(_03710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07972__A2 (.I(_03710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07971__A2 (.I(_03710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08004__A2 (.I(_03720_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08003__A2 (.I(_03720_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08002__A2 (.I(_03720_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08001__A2 (.I(_03720_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08000__A2 (.I(_03720_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07999__A2 (.I(_03720_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07998__A2 (.I(_03720_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07997__A2 (.I(_03720_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07996__A2 (.I(_03720_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07995__A2 (.I(_03720_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07994__A2 (.I(_03720_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07993__A2 (.I(_03720_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07992__A2 (.I(_03720_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07991__A2 (.I(_03720_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07990__A2 (.I(_03720_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07989__A2 (.I(_03720_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08022__A2 (.I(_03730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08021__A2 (.I(_03730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08020__A2 (.I(_03730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08019__A2 (.I(_03730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08018__A2 (.I(_03730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08017__A2 (.I(_03730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08016__A2 (.I(_03730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08015__A2 (.I(_03730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08014__A2 (.I(_03730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08013__A2 (.I(_03730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08012__A2 (.I(_03730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08011__A2 (.I(_03730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08010__A2 (.I(_03730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08009__A2 (.I(_03730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08008__A2 (.I(_03730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08007__A2 (.I(_03730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08040__A2 (.I(_03740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08039__A2 (.I(_03740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08038__A2 (.I(_03740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08037__A2 (.I(_03740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08036__A2 (.I(_03740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08035__A2 (.I(_03740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08034__A2 (.I(_03740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08033__A2 (.I(_03740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08032__A2 (.I(_03740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08031__A2 (.I(_03740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08030__A2 (.I(_03740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08029__A2 (.I(_03740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08028__A2 (.I(_03740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08027__A2 (.I(_03740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08026__A2 (.I(_03740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08025__A2 (.I(_03740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08058__A2 (.I(_03750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08057__A2 (.I(_03750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08056__A2 (.I(_03750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08055__A2 (.I(_03750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08054__A2 (.I(_03750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08053__A2 (.I(_03750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08052__A2 (.I(_03750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08051__A2 (.I(_03750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08050__A2 (.I(_03750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08049__A2 (.I(_03750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08048__A2 (.I(_03750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08047__A2 (.I(_03750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08046__A2 (.I(_03750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08045__A2 (.I(_03750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08044__A2 (.I(_03750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08043__A2 (.I(_03750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08076__A2 (.I(_03760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08075__A2 (.I(_03760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08074__A2 (.I(_03760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08073__A2 (.I(_03760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08072__A2 (.I(_03760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08071__A2 (.I(_03760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08070__A2 (.I(_03760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08069__A2 (.I(_03760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08068__A2 (.I(_03760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08067__A2 (.I(_03760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08066__A2 (.I(_03760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08065__A2 (.I(_03760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08064__A2 (.I(_03760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08063__A2 (.I(_03760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08062__A2 (.I(_03760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08061__A2 (.I(_03760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08094__A2 (.I(_03770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08093__A2 (.I(_03770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08092__A2 (.I(_03770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08091__A2 (.I(_03770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08090__A2 (.I(_03770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08089__A2 (.I(_03770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08088__A2 (.I(_03770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08087__A2 (.I(_03770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08086__A2 (.I(_03770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08085__A2 (.I(_03770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08084__A2 (.I(_03770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08083__A2 (.I(_03770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08082__A2 (.I(_03770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08081__A2 (.I(_03770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08080__A2 (.I(_03770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08079__A2 (.I(_03770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08112__A2 (.I(_03780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08111__A2 (.I(_03780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08110__A2 (.I(_03780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08109__A2 (.I(_03780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08108__A2 (.I(_03780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08107__A2 (.I(_03780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08106__A2 (.I(_03780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08105__A2 (.I(_03780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08104__A2 (.I(_03780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08103__A2 (.I(_03780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08102__A2 (.I(_03780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08101__A2 (.I(_03780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08100__A2 (.I(_03780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08099__A2 (.I(_03780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08098__A2 (.I(_03780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08097__A2 (.I(_03780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08130__A2 (.I(_03790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08129__A2 (.I(_03790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08128__A2 (.I(_03790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08127__A2 (.I(_03790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08126__A2 (.I(_03790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08125__A2 (.I(_03790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08124__A2 (.I(_03790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08123__A2 (.I(_03790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08122__A2 (.I(_03790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08121__A2 (.I(_03790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08120__A2 (.I(_03790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08119__A2 (.I(_03790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08118__A2 (.I(_03790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08117__A2 (.I(_03790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08116__A2 (.I(_03790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08115__A2 (.I(_03790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08231__A2 (.I(_03802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08164__A2 (.I(_03802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08160__B2 (.I(_03802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08152__A1 (.I(_03802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08145__A1 (.I(_03802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08140__A2 (.I(_03802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08136__A1 (.I(_03802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08242__A2 (.I(_03807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08240__A2 (.I(_03807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08237__A2 (.I(_03807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08232__A2 (.I(_03807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08229__A2 (.I(_03807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08226__A2 (.I(_03807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08223__A2 (.I(_03807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08220__A2 (.I(_03807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08217__A2 (.I(_03807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08214__A2 (.I(_03807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08160__C (.I(_03807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08157__I (.I(_03807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08141__A2 (.I(_03807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08140__A1 (.I(_03807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08242__B1 (.I(_03808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08239__A2 (.I(_03808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08236__A2 (.I(_03808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08232__B1 (.I(_03808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08229__B1 (.I(_03808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08225__A2 (.I(_03808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08222__A2 (.I(_03808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08219__A2 (.I(_03808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08216__A2 (.I(_03808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08213__A2 (.I(_03808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08173__I (.I(_03808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08171__A2 (.I(_03808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08167__B1 (.I(_03808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08141__B1 (.I(_03808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08211__A2 (.I(_03822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08208__A2 (.I(_03822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08205__A2 (.I(_03822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08202__A2 (.I(_03822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08199__A2 (.I(_03822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08196__A2 (.I(_03822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08193__A2 (.I(_03822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08190__A2 (.I(_03822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08187__A2 (.I(_03822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08184__A2 (.I(_03822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08181__A2 (.I(_03822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08178__A2 (.I(_03822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08175__A2 (.I(_03822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08169__A2 (.I(_03822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08167__A2 (.I(_03822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08161__A2 (.I(_03822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08240__B1 (.I(_03829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08237__B1 (.I(_03829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08226__B1 (.I(_03829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08223__B1 (.I(_03829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08220__B1 (.I(_03829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08217__B1 (.I(_03829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08214__B1 (.I(_03829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08170__I (.I(_03829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08166__C (.I(_03829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08245__B1 (.I(_03833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08228__A2 (.I(_03833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08211__B1 (.I(_03833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08208__B1 (.I(_03833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08205__B1 (.I(_03833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08202__B1 (.I(_03833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08199__B1 (.I(_03833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08196__B1 (.I(_03833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08193__B1 (.I(_03833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08190__B1 (.I(_03833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08187__B1 (.I(_03833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08184__B1 (.I(_03833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08181__B1 (.I(_03833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08178__B1 (.I(_03833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08175__B1 (.I(_03833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08171__B1 (.I(_03833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08247__A2 (.I(_03835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08245__A2 (.I(_03835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08235__A2 (.I(_03835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08210__A2 (.I(_03835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08207__A2 (.I(_03835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08204__A2 (.I(_03835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08201__A2 (.I(_03835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08198__A2 (.I(_03835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08195__A2 (.I(_03835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08192__A2 (.I(_03835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08189__A2 (.I(_03835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08186__A2 (.I(_03835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08183__A2 (.I(_03835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08180__A2 (.I(_03835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08177__A2 (.I(_03835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08174__A2 (.I(_03835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08246__B1 (.I(_03874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08243__A2 (.I(_03874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08234__B1 (.I(_03874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08233__A2 (.I(_03874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08265__A2 (.I(_03885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08264__A2 (.I(_03885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08263__A2 (.I(_03885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08262__A2 (.I(_03885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08261__A2 (.I(_03885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08260__A2 (.I(_03885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08259__A2 (.I(_03885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08258__A2 (.I(_03885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08257__A2 (.I(_03885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08256__A2 (.I(_03885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08255__A2 (.I(_03885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08254__A2 (.I(_03885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08253__A2 (.I(_03885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08252__A2 (.I(_03885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08251__A2 (.I(_03885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08250__A2 (.I(_03885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08389__A1 (.I(_03895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08268__I (.I(_03895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09690__A1 (.I(_03896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08948__A1 (.I(_03896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08644__C (.I(_03896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08639__B (.I(_03896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08629__A1 (.I(_03896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08606__C (.I(_03896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08564__B (.I(_03896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08562__A1 (.I(_03896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08524__A1 (.I(_03896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08504__A1 (.I(_03896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08478__C (.I(_03896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08468__B (.I(_03896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08461__A1 (.I(_03896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08356__C (.I(_03896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08327__C (.I(_03896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08269__I (.I(_03896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09524__A2 (.I(_03897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09045__A2 (.I(_03897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08963__A2 (.I(_03897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08953__B (.I(_03897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08939__B2 (.I(_03897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08928__A2 (.I(_03897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08645__A2 (.I(_03897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08592__A2 (.I(_03897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08579__A2 (.I(_03897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08576__A2 (.I(_03897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08573__A2 (.I(_03897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08570__A2 (.I(_03897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08566__B2 (.I(_03897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08328__A2 (.I(_03897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08326__A1 (.I(_03897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08325__A2 (.I(_03897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08560__A1 (.I(_03899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08491__B (.I(_03899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08454__A1 (.I(_03899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08395__A1 (.I(_03899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08392__A1 (.I(_03899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08391__B2 (.I(_03899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08366__A1 (.I(_03899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08324__A1 (.I(_03899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08318__A4 (.I(_03899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08959__A1 (.I(_03901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08509__A1 (.I(_03901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08493__A1 (.I(_03901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08455__B2 (.I(_03901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08407__A1 (.I(_03901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08404__A1 (.I(_03901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08394__A1 (.I(_03901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08344__A1 (.I(_03901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08341__A1 (.I(_03901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08311__A1 (.I(_03901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08282__A1 (.I(_03901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08276__A1 (.I(_03901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08954__A1 (.I(_03903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08558__A1 (.I(_03903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08494__B1 (.I(_03903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08363__A2 (.I(_03903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08287__A2 (.I(_03903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08282__A2 (.I(_03903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08276__A2 (.I(_03903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08591__A2 (.I(_03904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08397__A2 (.I(_03904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08386__A2 (.I(_03904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08338__A1 (.I(_03904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08284__A1 (.I(_03904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08617__A2 (.I(_03906_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08596__A2 (.I(_03906_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08586__A2 (.I(_03906_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08534__A1 (.I(_03906_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08475__A1 (.I(_03906_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08442__A1 (.I(_03906_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08337__A1 (.I(_03906_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08336__A1 (.I(_03906_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08335__A2 (.I(_03906_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08321__A1 (.I(_03906_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08291__A1 (.I(_03906_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08290__A1 (.I(_03906_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08281__A1 (.I(_03906_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08934__A2 (.I(_03908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08588__A1 (.I(_03908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08585__A3 (.I(_03908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08560__A2 (.I(_03908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08554__B2 (.I(_03908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08533__A1 (.I(_03908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08485__A2 (.I(_03908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08474__A2 (.I(_03908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08414__A2 (.I(_03908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08365__A2 (.I(_03908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08362__A2 (.I(_03908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08356__A2 (.I(_03908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08291__A2 (.I(_03908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08281__A2 (.I(_03908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08934__B1 (.I(_03909_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08617__B1 (.I(_03909_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08595__A1 (.I(_03909_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08560__B1 (.I(_03909_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08513__B2 (.I(_03909_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08485__B1 (.I(_03909_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08414__B1 (.I(_03909_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08345__A1 (.I(_03909_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08283__A1 (.I(_03909_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08946__A2 (.I(_03910_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08935__B2 (.I(_03910_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08933__A1 (.I(_03910_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08626__A2 (.I(_03910_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08623__B (.I(_03910_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08584__A1 (.I(_03910_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08533__C (.I(_03910_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08522__A2 (.I(_03910_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08514__B2 (.I(_03910_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08457__A1 (.I(_03910_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08409__A1 (.I(_03910_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08396__A1 (.I(_03910_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08283__A2 (.I(_03910_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08636__B (.I(_03912_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08606__A1 (.I(_03912_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08605__B (.I(_03912_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08562__A2 (.I(_03912_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08478__A1 (.I(_03912_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08477__C (.I(_03912_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08361__B (.I(_03912_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08356__B1 (.I(_03912_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08333__A2 (.I(_03912_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08327__A2 (.I(_03912_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08324__A2 (.I(_03912_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08559__B2 (.I(_03914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08494__A2 (.I(_03914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08486__A1 (.I(_03914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08413__A1 (.I(_03914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08363__A1 (.I(_03914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08356__A1 (.I(_03914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08335__A1 (.I(_03914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08287__A1 (.I(_03914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08625__C (.I(_03915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08587__B (.I(_03915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08444__B (.I(_03915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08416__B (.I(_03915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08368__A1 (.I(_03915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08361__A1 (.I(_03915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08327__B1 (.I(_03915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08324__B1 (.I(_03915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08490__A3 (.I(_03917_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08443__A1 (.I(_03917_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08392__A2 (.I(_03917_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08345__A2 (.I(_03917_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08337__A2 (.I(_03917_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08302__A1 (.I(_03917_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08290__A2 (.I(_03917_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08954__A2 (.I(_03918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08624__A1 (.I(_03918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08588__A2 (.I(_03918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08581__A2 (.I(_03918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08541__A2 (.I(_03918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08528__A2 (.I(_03918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08518__A2 (.I(_03918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08483__A2 (.I(_03918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08451__A2 (.I(_03918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08385__A2 (.I(_03918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08379__A2 (.I(_03918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08361__A2 (.I(_03918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08327__B2 (.I(_03918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08303__A1 (.I(_03918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08962__A2 (.I(_03922_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08638__A1 (.I(_03922_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08633__A1 (.I(_03922_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08540__A1 (.I(_03922_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08539__B (.I(_03922_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08485__A1 (.I(_03922_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08483__A1 (.I(_03922_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08446__A1 (.I(_03922_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08377__C (.I(_03922_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08346__A1 (.I(_03922_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08298__A1 (.I(_03922_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08955__B (.I(_03923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08625__A1 (.I(_03923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08623__A1 (.I(_03923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08540__A2 (.I(_03923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08539__A1 (.I(_03923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08528__A1 (.I(_03923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08346__A2 (.I(_03923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08298__A2 (.I(_03923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08943__A1 (.I(_03924_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08942__A1 (.I(_03924_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08617__A1 (.I(_03924_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08614__B (.I(_03924_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08587__A1 (.I(_03924_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08522__A1 (.I(_03924_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08518__A1 (.I(_03924_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08298__A3 (.I(_03924_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08589__B (.I(_03925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08563__A1 (.I(_03925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08560__B2 (.I(_03925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08557__A1 (.I(_03925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08554__A1 (.I(_03925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08553__A1 (.I(_03925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08551__A1 (.I(_03925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08456__C2 (.I(_03925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08454__B2 (.I(_03925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08451__A1 (.I(_03925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08298__A4 (.I(_03925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08932__A1 (.I(_03928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08602__A1 (.I(_03928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08601__A1 (.I(_03928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08490__A2 (.I(_03928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08351__A2 (.I(_03928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08301__A2 (.I(_03928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08598__A2 (.I(_03929_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08519__A2 (.I(_03929_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08450__A2 (.I(_03929_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08449__A2 (.I(_03929_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08302__A3 (.I(_03929_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08939__A1 (.I(_03932_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08934__B2 (.I(_03932_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08931__A1 (.I(_03932_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08930__A1 (.I(_03932_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08599__A1 (.I(_03932_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08596__A1 (.I(_03932_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08541__A1 (.I(_03932_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08513__A1 (.I(_03932_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08510__A1 (.I(_03932_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08305__A2 (.I(_03932_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08555__A1 (.I(_03935_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08539__A2 (.I(_03935_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08529__A1 (.I(_03935_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08494__A1 (.I(_03935_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08445__A1 (.I(_03935_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08415__A1 (.I(_03935_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08369__A1 (.I(_03935_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08308__A2 (.I(_03935_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08391__A1 (.I(_03936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08334__A1 (.I(_03936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08323__A1 (.I(_03936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08511__B (.I(_03938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08486__B (.I(_03938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08454__C (.I(_03938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08413__A2 (.I(_03938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08408__A1 (.I(_03938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08406__B (.I(_03938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08391__C (.I(_03938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08344__A2 (.I(_03938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08334__A2 (.I(_03938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08311__A2 (.I(_03938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08946__A1 (.I(_03940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08598__A1 (.I(_03940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08508__A1 (.I(_03940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08486__A2 (.I(_03940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08483__B2 (.I(_03940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08414__A1 (.I(_03940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08377__A2 (.I(_03940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08364__A1 (.I(_03940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08359__B1 (.I(_03940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08314__A1 (.I(_03940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08476__A1 (.I(_03941_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08473__A1 (.I(_03941_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08456__A2 (.I(_03941_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08451__B2 (.I(_03941_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08364__A2 (.I(_03941_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08314__A2 (.I(_03941_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08934__A1 (.I(_03944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08931__B2 (.I(_03944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08511__A1 (.I(_03944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08507__A1 (.I(_03944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08408__B2 (.I(_03944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08402__A1 (.I(_03944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08379__B2 (.I(_03944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08327__A1 (.I(_03944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08318__A2 (.I(_03944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08944__A1 (.I(_03945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08414__C2 (.I(_03945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08385__B2 (.I(_03945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08318__A3 (.I(_03945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08956__A1 (.I(_03947_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08947__A2 (.I(_03947_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08591__A1 (.I(_03947_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08476__B2 (.I(_03947_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08442__A2 (.I(_03947_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08405__A1 (.I(_03947_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08375__A2 (.I(_03947_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08350__A2 (.I(_03947_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08336__A2 (.I(_03947_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08320__A2 (.I(_03947_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08960__B (.I(_03948_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08930__A3 (.I(_03948_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08557__A2 (.I(_03948_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08334__A3 (.I(_03948_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08321__A2 (.I(_03948_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08360__A1 (.I(_03950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08323__A2 (.I(_03950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08328__B (.I(_03954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08950__C (.I(_03955_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08927__A1 (.I(_03955_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08637__A1 (.I(_03955_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08630__A2 (.I(_03955_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08619__A2 (.I(_03955_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08607__A2 (.I(_03955_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08591__C (.I(_03955_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08543__B2 (.I(_03955_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08501__A1 (.I(_03955_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08499__A1 (.I(_03955_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08479__A2 (.I(_03955_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08462__A1 (.I(_03955_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08421__C (.I(_03955_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08410__B2 (.I(_03955_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08381__C (.I(_03955_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08330__I (.I(_03955_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08962__A1 (.I(_03956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08957__A1 (.I(_03956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08936__A1 (.I(_03956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08500__A2 (.I(_03956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08459__A2 (.I(_03956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08422__A2 (.I(_03956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08411__A2 (.I(_03956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08400__A2 (.I(_03956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08388__A2 (.I(_03956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08387__A1 (.I(_03956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08382__A2 (.I(_03956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08371__A2 (.I(_03956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08370__A1 (.I(_03956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08359__A2 (.I(_03956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08358__A2 (.I(_03956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08343__A2 (.I(_03956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08947__A1 (.I(_03958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08519__A1 (.I(_03958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08418__B (.I(_03958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08343__B1 (.I(_03958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08621__A1 (.I(_03959_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08536__C2 (.I(_03959_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08526__C2 (.I(_03959_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08500__B1 (.I(_03959_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08359__B2 (.I(_03959_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08343__B2 (.I(_03959_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08603__A2 (.I(_03961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08494__B2 (.I(_03961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08372__A2 (.I(_03961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08342__A2 (.I(_03961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08961__A2 (.I(_03962_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08947__B1 (.I(_03962_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08930__A4 (.I(_03962_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08557__A3 (.I(_03962_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08555__A2 (.I(_03962_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08392__A3 (.I(_03962_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08337__B (.I(_03962_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08508__A2 (.I(_03963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08491__A1 (.I(_03963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08352__I (.I(_03963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08341__A2 (.I(_03963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08961__A1 (.I(_03965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08941__B (.I(_03965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08933__B (.I(_03965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08628__B (.I(_03965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08590__A1 (.I(_03965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08421__A1 (.I(_03965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08420__C (.I(_03965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08389__A2 (.I(_03965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08381__A1 (.I(_03965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08372__A1 (.I(_03965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08340__A2 (.I(_03965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09525__A1 (.I(_03966_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08535__A1 (.I(_03966_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08523__A1 (.I(_03966_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08514__C (.I(_03966_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08495__B (.I(_03966_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08487__A1 (.I(_03966_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08457__B (.I(_03966_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08341__B (.I(_03966_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08956__B1 (.I(_03969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08932__C (.I(_03969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08634__B (.I(_03969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08601__C (.I(_03969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08552__A1 (.I(_03969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08418__A1 (.I(_03969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08386__B1 (.I(_03969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08380__B (.I(_03969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08357__A1 (.I(_03969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08598__C (.I(_03972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08597__A1 (.I(_03972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08449__C (.I(_03972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08405__A2 (.I(_03972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08381__A2 (.I(_03972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08376__A2 (.I(_03972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08366__B2 (.I(_03972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08351__B (.I(_03972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08626__A1 (.I(_03974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08553__A2 (.I(_03974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08529__A2 (.I(_03974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08456__A1 (.I(_03974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08445__A2 (.I(_03974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08416__A1 (.I(_03974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08406__A1 (.I(_03974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08386__A1 (.I(_03974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08375__A1 (.I(_03974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08365__A1 (.I(_03974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08362__A1 (.I(_03974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08350__A1 (.I(_03974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08931__A2 (.I(_03975_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08624__A2 (.I(_03975_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08598__B (.I(_03975_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08511__A2 (.I(_03975_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08507__A2 (.I(_03975_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08454__A2 (.I(_03975_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08449__B (.I(_03975_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08407__A2 (.I(_03975_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08351__C (.I(_03975_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08358__B (.I(_03982_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08943__A3 (.I(_03985_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08597__A2 (.I(_03985_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08584__A2 (.I(_03985_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08456__C1 (.I(_03985_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08369__B1 (.I(_03985_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08941__A1 (.I(_03986_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08602__A2 (.I(_03986_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08586__A1 (.I(_03986_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08417__A1 (.I(_03986_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08369__B2 (.I(_03986_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08944__A2 (.I(_03988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08931__B1 (.I(_03988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08518__B1 (.I(_03988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08510__A2 (.I(_03988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08454__B1 (.I(_03988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08451__B1 (.I(_03988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08414__C1 (.I(_03988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08402__A2 (.I(_03988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08395__A2 (.I(_03988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08366__B1 (.I(_03988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08574__B2 (.I(_03993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08371__B (.I(_03993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08599__A2 (.I(_03998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08554__A2 (.I(_03998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08540__C (.I(_03998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08446__A4 (.I(_03998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08377__B (.I(_03998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08585__A1 (.I(_04000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08581__A1 (.I(_04000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08556__A2 (.I(_04000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08518__B2 (.I(_04000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08492__A1 (.I(_04000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08449__A1 (.I(_04000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08446__A3 (.I(_04000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08444__A1 (.I(_04000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08403__A1 (.I(_04000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08393__A1 (.I(_04000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08385__A1 (.I(_04000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08379__A1 (.I(_04000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08577__B2 (.I(_04003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08382__B (.I(_04003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08540__B1 (.I(_04004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08384__A2 (.I(_04004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08580__B2 (.I(_04008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08388__B (.I(_04008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08939__A2 (.I(_04009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08645__B1 (.I(_04009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08563__A2 (.I(_04009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08543__A1 (.I(_04009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08516__C2 (.I(_04009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08488__C2 (.I(_04009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08458__A1 (.I(_04009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08410__A1 (.I(_04009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08399__A1 (.I(_04009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08399__A2 (.I(_04010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08634__A1 (.I(_04013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08624__B (.I(_04013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08613__A1 (.I(_04013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08394__A3 (.I(_04013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08571__B2 (.I(_04019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08464__A1 (.I(_04019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08400__B (.I(_04019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08410__A2 (.I(_04020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08960__A1 (.I(_04024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08492__A2 (.I(_04024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08447__A1 (.I(_04024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08416__A3 (.I(_04024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08406__A2 (.I(_04024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08466__A1 (.I(_04029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08411__B (.I(_04029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08421__A2 (.I(_04030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08414__B2 (.I(_04030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08960__C (.I(_04031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08956__A2 (.I(_04031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08954__B (.I(_04031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08947__A3 (.I(_04031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08617__C (.I(_04031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08615__A1 (.I(_04031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08603__A1 (.I(_04031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08596__B (.I(_04031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08560__C (.I(_04031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08485__C (.I(_04031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08477__A1 (.I(_04031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08476__C (.I(_04031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08420__A1 (.I(_04031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08469__B2 (.I(_04039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08422__B (.I(_04039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08440__A2 (.I(_04041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08439__A2 (.I(_04041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08438__A2 (.I(_04041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08437__A2 (.I(_04041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08436__A2 (.I(_04041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08435__A2 (.I(_04041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08434__A2 (.I(_04041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08433__A2 (.I(_04041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08432__A2 (.I(_04041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08431__A2 (.I(_04041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08430__A2 (.I(_04041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08429__A2 (.I(_04041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08428__A2 (.I(_04041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08427__A2 (.I(_04041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08426__A2 (.I(_04041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08425__A2 (.I(_04041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08458__A2 (.I(_04050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08456__B2 (.I(_04050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08596__C (.I(_04051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08522__A3 (.I(_04051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08513__A2 (.I(_04051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08476__A2 (.I(_04051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08443__A2 (.I(_04051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08625__A2 (.I(_04052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08613__A2 (.I(_04052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08600__A2 (.I(_04052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08587__A2 (.I(_04052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08582__C (.I(_04052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08551__A2 (.I(_04052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08529__B (.I(_04052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08448__A1 (.I(_04052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08444__A2 (.I(_04052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08506__A1 (.I(_04067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08459__B (.I(_04067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08468__A2 (.I(_04068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08462__A2 (.I(_04068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08461__A2 (.I(_04068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08488__A2 (.I(_04069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08481__A1 (.I(_04069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08480__A2 (.I(_04069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08469__A2 (.I(_04069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08465__A2 (.I(_04069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08463__A2 (.I(_04069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08488__B1 (.I(_04070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08465__B1 (.I(_04070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08463__B1 (.I(_04070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08478__A2 (.I(_04075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08476__B1 (.I(_04075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08481__A2 (.I(_04083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08488__C1 (.I(_04088_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08485__B2 (.I(_04088_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08507__A3 (.I(_04093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08491__A2 (.I(_04093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08495__A2 (.I(_04097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08500__B2 (.I(_04099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08524__A2 (.I(_04101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08504__A2 (.I(_04101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08501__A2 (.I(_04101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08499__A2 (.I(_04101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08549__B (.I(_04106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08516__B1 (.I(_04106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08505__B1 (.I(_04106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08600__A3 (.I(_04111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08514__A1 (.I(_04111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08516__C1 (.I(_04113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08513__B1 (.I(_04113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08523__A2 (.I(_04121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08536__C1 (.I(_04131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08533__A2 (.I(_04131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09046__A1 (.I(_04141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08550__A1 (.I(_04141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08929__B2 (.I(_04160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08566__A1 (.I(_04160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08620__A1 (.I(_04164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08579__B (.I(_04164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08569__I (.I(_04164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08642__A1 (.I(_04165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08641__A2 (.I(_04165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08632__A1 (.I(_04165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08631__A2 (.I(_04165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08610__A2 (.I(_04165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08609__A1 (.I(_04165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08608__A2 (.I(_04165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08593__A2 (.I(_04165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08592__B (.I(_04165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08580__A2 (.I(_04165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08577__A2 (.I(_04165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08576__B (.I(_04165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08574__A2 (.I(_04165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08573__B (.I(_04165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08571__A2 (.I(_04165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08570__B (.I(_04165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08593__B1 (.I(_04183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08609__A2 (.I(_04197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08621__A2 (.I(_04202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08617__B2 (.I(_04202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08632__A2 (.I(_04218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08642__A3 (.I(_04228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08645__C (.I(_04231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08668__A2 (.I(_04237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08667__A2 (.I(_04237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08666__A2 (.I(_04237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08665__A2 (.I(_04237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08664__A2 (.I(_04237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08663__A2 (.I(_04237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08662__A2 (.I(_04237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08661__A2 (.I(_04237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08660__A2 (.I(_04237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08659__A2 (.I(_04237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08658__A2 (.I(_04237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08657__A2 (.I(_04237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08656__A2 (.I(_04237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08655__A2 (.I(_04237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08654__A2 (.I(_04237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08653__A2 (.I(_04237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08686__A2 (.I(_04247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08685__A2 (.I(_04247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08684__A2 (.I(_04247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08683__A2 (.I(_04247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08682__A2 (.I(_04247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08681__A2 (.I(_04247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08680__A2 (.I(_04247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08679__A2 (.I(_04247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08678__A2 (.I(_04247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08677__A2 (.I(_04247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08676__A2 (.I(_04247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08675__A2 (.I(_04247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08674__A2 (.I(_04247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08673__A2 (.I(_04247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08672__A2 (.I(_04247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08671__A2 (.I(_04247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08720__S (.I(_04257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08718__S (.I(_04257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08716__S (.I(_04257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08714__S (.I(_04257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08712__S (.I(_04257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08710__S (.I(_04257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08708__S (.I(_04257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08706__S (.I(_04257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08704__S (.I(_04257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08702__S (.I(_04257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08700__S (.I(_04257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08698__S (.I(_04257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08696__S (.I(_04257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08694__S (.I(_04257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08692__S (.I(_04257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08690__S (.I(_04257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08759__A1 (.I(_04288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08751__A1 (.I(_04288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08760__S (.I(_04293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08757__A2 (.I(_04293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08756__A2 (.I(_04293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08779__A2 (.I(_04299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08778__A2 (.I(_04299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08777__A2 (.I(_04299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08776__A2 (.I(_04299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08775__A2 (.I(_04299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08774__A2 (.I(_04299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08773__A2 (.I(_04299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08772__A2 (.I(_04299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08771__A2 (.I(_04299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08770__A2 (.I(_04299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08769__A2 (.I(_04299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08768__A2 (.I(_04299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08767__A2 (.I(_04299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08766__A2 (.I(_04299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08765__A2 (.I(_04299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08764__A2 (.I(_04299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09692__A1 (.I(_04309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08812__A2 (.I(_04309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08810__A2 (.I(_04309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08808__A2 (.I(_04309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08806__A2 (.I(_04309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08804__A2 (.I(_04309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08802__A2 (.I(_04309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08800__A2 (.I(_04309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08798__A2 (.I(_04309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08796__A2 (.I(_04309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08794__A2 (.I(_04309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08792__A2 (.I(_04309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08790__A2 (.I(_04309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08788__A2 (.I(_04309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08786__A2 (.I(_04309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08784__A2 (.I(_04309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08815__B1 (.I(_04311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08812__B1 (.I(_04311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08810__B1 (.I(_04311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08808__B1 (.I(_04311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08806__B1 (.I(_04311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08804__B1 (.I(_04311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08802__B1 (.I(_04311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08800__B1 (.I(_04311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08798__B1 (.I(_04311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08796__B1 (.I(_04311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08794__B1 (.I(_04311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08792__B1 (.I(_04311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08790__B1 (.I(_04311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08788__B1 (.I(_04311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08786__B1 (.I(_04311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08784__B1 (.I(_04311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08846__A2 (.I(_04327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08844__A2 (.I(_04327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08842__A2 (.I(_04327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08840__A2 (.I(_04327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08838__A2 (.I(_04327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08836__A2 (.I(_04327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08834__A2 (.I(_04327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08832__A2 (.I(_04327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08830__A2 (.I(_04327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08828__A2 (.I(_04327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08826__A2 (.I(_04327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08824__A2 (.I(_04327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08822__A2 (.I(_04327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08820__A2 (.I(_04327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08818__A2 (.I(_04327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08815__A2 (.I(_04327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08851__B1 (.I(_04329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08846__B1 (.I(_04329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08844__B1 (.I(_04329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08842__B1 (.I(_04329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08840__B1 (.I(_04329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08838__B1 (.I(_04329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08836__B1 (.I(_04329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08834__B1 (.I(_04329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08832__B1 (.I(_04329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08830__B1 (.I(_04329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08828__B1 (.I(_04329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08826__B1 (.I(_04329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08824__B1 (.I(_04329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08822__B1 (.I(_04329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08820__B1 (.I(_04329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08818__B1 (.I(_04329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08851__B2 (.I(_04347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09636__A2 (.I(_04349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09618__A2 (.I(_04349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09433__A2 (.I(_04349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09397__A2 (.I(_04349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09281__A2 (.I(_04349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09245__A2 (.I(_04349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09227__A2 (.I(_04349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09209__A2 (.I(_04349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09173__A2 (.I(_04349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09155__A2 (.I(_04349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09137__A2 (.I(_04349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09119__A2 (.I(_04349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09101__A2 (.I(_04349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09027__A2 (.I(_04349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08965__A2 (.I(_04349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08854__A2 (.I(_04349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08871__A2 (.I(_04351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08870__A2 (.I(_04351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08869__A2 (.I(_04351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08868__A2 (.I(_04351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08867__A2 (.I(_04351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08866__A2 (.I(_04351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08865__A2 (.I(_04351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08864__A2 (.I(_04351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08863__A2 (.I(_04351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08862__A2 (.I(_04351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08861__A2 (.I(_04351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08860__A2 (.I(_04351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08859__A2 (.I(_04351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08858__A2 (.I(_04351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08857__A2 (.I(_04351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08856__A2 (.I(_04351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08889__A2 (.I(_04361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08888__A2 (.I(_04361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08887__A2 (.I(_04361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08886__A2 (.I(_04361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08885__A2 (.I(_04361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08884__A2 (.I(_04361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08883__A2 (.I(_04361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08882__A2 (.I(_04361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08881__A2 (.I(_04361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08880__A2 (.I(_04361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08879__A2 (.I(_04361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08878__A2 (.I(_04361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08877__A2 (.I(_04361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08876__A2 (.I(_04361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08875__A2 (.I(_04361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08874__A2 (.I(_04361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08907__A2 (.I(_04371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08906__A2 (.I(_04371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08905__A2 (.I(_04371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08904__A2 (.I(_04371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08903__A2 (.I(_04371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08902__A2 (.I(_04371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08901__A2 (.I(_04371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08900__A2 (.I(_04371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08899__A2 (.I(_04371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08898__A2 (.I(_04371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08897__A2 (.I(_04371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08896__A2 (.I(_04371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08895__A2 (.I(_04371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08894__A2 (.I(_04371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08893__A2 (.I(_04371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08892__A2 (.I(_04371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08925__A2 (.I(_04381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08924__A2 (.I(_04381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08923__A2 (.I(_04381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08922__A2 (.I(_04381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08921__A2 (.I(_04381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08920__A2 (.I(_04381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08919__A2 (.I(_04381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08918__A2 (.I(_04381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08917__A2 (.I(_04381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08916__A2 (.I(_04381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08915__A2 (.I(_04381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08914__A2 (.I(_04381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08913__A2 (.I(_04381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08912__A2 (.I(_04381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08911__A2 (.I(_04381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08910__A2 (.I(_04381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08957__A2 (.I(_04417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08982__A2 (.I(_04425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08981__A2 (.I(_04425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08980__A2 (.I(_04425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08979__A2 (.I(_04425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08978__A2 (.I(_04425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08977__A2 (.I(_04425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08976__A2 (.I(_04425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08975__A2 (.I(_04425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08974__A2 (.I(_04425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08973__A2 (.I(_04425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08972__A2 (.I(_04425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08971__A2 (.I(_04425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08970__A2 (.I(_04425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08969__A2 (.I(_04425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08968__A2 (.I(_04425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08967__A2 (.I(_04425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09302__A1 (.I(_04434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09284__A1 (.I(_04434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09266__A1 (.I(_04434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09248__A1 (.I(_04434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09230__A1 (.I(_04434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09212__A1 (.I(_04434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09194__A1 (.I(_04434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09176__A1 (.I(_04434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09158__A1 (.I(_04434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09140__A1 (.I(_04434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09122__A1 (.I(_04434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09104__A1 (.I(_04434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09053__A1 (.I(_04434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09030__A1 (.I(_04434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09012__A1 (.I(_04434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08987__A1 (.I(_04434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09008__A2 (.I(_04436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09007__A2 (.I(_04436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09005__A2 (.I(_04436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09004__A2 (.I(_04436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09002__A2 (.I(_04436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09001__A2 (.I(_04436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08999__A2 (.I(_04436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08998__A2 (.I(_04436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08996__A2 (.I(_04436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08995__A2 (.I(_04436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08993__A2 (.I(_04436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08992__A2 (.I(_04436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08990__A2 (.I(_04436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08989__A2 (.I(_04436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08987__A2 (.I(_04436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08986__A2 (.I(_04436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09304__A1 (.I(_04438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09286__A1 (.I(_04438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09268__A1 (.I(_04438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09250__A1 (.I(_04438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09232__A1 (.I(_04438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09214__A1 (.I(_04438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09196__A1 (.I(_04438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09178__A1 (.I(_04438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09160__A1 (.I(_04438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09142__A1 (.I(_04438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09124__A1 (.I(_04438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09106__A1 (.I(_04438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09055__A1 (.I(_04438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09032__A1 (.I(_04438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09014__A1 (.I(_04438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08990__A1 (.I(_04438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09306__A1 (.I(_04440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09288__A1 (.I(_04440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09270__A1 (.I(_04440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09252__A1 (.I(_04440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09234__A1 (.I(_04440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09216__A1 (.I(_04440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09198__A1 (.I(_04440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09180__A1 (.I(_04440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09162__A1 (.I(_04440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09144__A1 (.I(_04440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09126__A1 (.I(_04440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09108__A1 (.I(_04440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09057__A1 (.I(_04440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09034__A1 (.I(_04440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09016__A1 (.I(_04440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08993__A1 (.I(_04440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09308__A1 (.I(_04442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09290__A1 (.I(_04442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09272__A1 (.I(_04442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09254__A1 (.I(_04442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09236__A1 (.I(_04442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09218__A1 (.I(_04442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09200__A1 (.I(_04442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09182__A1 (.I(_04442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09164__A1 (.I(_04442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09146__A1 (.I(_04442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09128__A1 (.I(_04442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09110__A1 (.I(_04442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09059__A1 (.I(_04442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09036__A1 (.I(_04442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09018__A1 (.I(_04442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08996__A1 (.I(_04442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09310__A1 (.I(_04444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09292__A1 (.I(_04444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09274__A1 (.I(_04444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09256__A1 (.I(_04444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09238__A1 (.I(_04444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09220__A1 (.I(_04444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09202__A1 (.I(_04444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09184__A1 (.I(_04444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09166__A1 (.I(_04444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09148__A1 (.I(_04444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09130__A1 (.I(_04444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09112__A1 (.I(_04444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09061__A1 (.I(_04444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09038__A1 (.I(_04444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09020__A1 (.I(_04444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08999__A1 (.I(_04444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09312__A1 (.I(_04446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09294__A1 (.I(_04446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09276__A1 (.I(_04446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09258__A1 (.I(_04446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09240__A1 (.I(_04446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09222__A1 (.I(_04446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09204__A1 (.I(_04446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09186__A1 (.I(_04446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09168__A1 (.I(_04446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09150__A1 (.I(_04446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09132__A1 (.I(_04446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09114__A1 (.I(_04446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09063__A1 (.I(_04446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09040__A1 (.I(_04446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09022__A1 (.I(_04446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09002__A1 (.I(_04446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09314__A1 (.I(_04448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09296__A1 (.I(_04448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09278__A1 (.I(_04448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09260__A1 (.I(_04448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09242__A1 (.I(_04448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09224__A1 (.I(_04448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09206__A1 (.I(_04448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09188__A1 (.I(_04448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09170__A1 (.I(_04448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09152__A1 (.I(_04448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09134__A1 (.I(_04448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09116__A1 (.I(_04448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09065__A1 (.I(_04448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09042__A1 (.I(_04448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09024__A1 (.I(_04448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09005__A1 (.I(_04448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09316__A1 (.I(_04450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09298__A1 (.I(_04450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09280__A1 (.I(_04450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09262__A1 (.I(_04450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09244__A1 (.I(_04450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09226__A1 (.I(_04450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09208__A1 (.I(_04450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09190__A1 (.I(_04450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09172__A1 (.I(_04450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09154__A1 (.I(_04450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09136__A1 (.I(_04450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09118__A1 (.I(_04450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09067__A1 (.I(_04450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09044__A1 (.I(_04450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09026__A1 (.I(_04450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09008__A1 (.I(_04450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09026__A2 (.I(_04453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09025__A2 (.I(_04453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09024__A2 (.I(_04453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09023__A2 (.I(_04453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09022__A2 (.I(_04453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09021__A2 (.I(_04453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09020__A2 (.I(_04453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09019__A2 (.I(_04453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09018__A2 (.I(_04453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09017__A2 (.I(_04453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09016__A2 (.I(_04453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09015__A2 (.I(_04453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09014__A2 (.I(_04453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09013__A2 (.I(_04453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09012__A2 (.I(_04453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09011__A2 (.I(_04453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09044__A2 (.I(_04463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09043__A2 (.I(_04463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09042__A2 (.I(_04463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09041__A2 (.I(_04463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09040__A2 (.I(_04463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09039__A2 (.I(_04463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09038__A2 (.I(_04463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09037__A2 (.I(_04463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09036__A2 (.I(_04463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09035__A2 (.I(_04463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09034__A2 (.I(_04463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09033__A2 (.I(_04463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09032__A2 (.I(_04463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09031__A2 (.I(_04463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09030__A2 (.I(_04463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09029__A2 (.I(_04463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09067__A2 (.I(_04476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09066__A2 (.I(_04476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09065__A2 (.I(_04476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09064__A2 (.I(_04476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09063__A2 (.I(_04476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09062__A2 (.I(_04476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09061__A2 (.I(_04476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09060__A2 (.I(_04476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09059__A2 (.I(_04476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09058__A2 (.I(_04476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09057__A2 (.I(_04476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09056__A2 (.I(_04476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09055__A2 (.I(_04476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09054__A2 (.I(_04476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09053__A2 (.I(_04476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09052__A2 (.I(_04476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09097__S (.I(_04485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09095__S (.I(_04485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09093__S (.I(_04485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09092__A2 (.I(_04485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09091__A2 (.I(_04485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09089__S (.I(_04485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09087__S (.I(_04485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09085__S (.I(_04485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09083__S (.I(_04485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09081__S (.I(_04485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09079__S (.I(_04485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09077__S (.I(_04485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09075__S (.I(_04485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09073__S (.I(_04485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09071__S (.I(_04485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09069__S (.I(_04485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09118__A2 (.I(_04503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09117__A2 (.I(_04503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09116__A2 (.I(_04503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09115__A2 (.I(_04503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09114__A2 (.I(_04503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09113__A2 (.I(_04503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09112__A2 (.I(_04503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09111__A2 (.I(_04503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09110__A2 (.I(_04503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09109__A2 (.I(_04503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09108__A2 (.I(_04503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09107__A2 (.I(_04503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09106__A2 (.I(_04503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09105__A2 (.I(_04503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09104__A2 (.I(_04503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09103__A2 (.I(_04503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09136__A2 (.I(_04513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09135__A2 (.I(_04513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09134__A2 (.I(_04513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09133__A2 (.I(_04513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09132__A2 (.I(_04513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09131__A2 (.I(_04513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09130__A2 (.I(_04513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09129__A2 (.I(_04513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09128__A2 (.I(_04513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09127__A2 (.I(_04513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09126__A2 (.I(_04513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09125__A2 (.I(_04513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09124__A2 (.I(_04513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09123__A2 (.I(_04513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09122__A2 (.I(_04513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09121__A2 (.I(_04513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09154__A2 (.I(_04523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09153__A2 (.I(_04523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09152__A2 (.I(_04523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09151__A2 (.I(_04523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09150__A2 (.I(_04523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09149__A2 (.I(_04523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09148__A2 (.I(_04523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09147__A2 (.I(_04523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09146__A2 (.I(_04523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09145__A2 (.I(_04523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09144__A2 (.I(_04523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09143__A2 (.I(_04523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09142__A2 (.I(_04523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09141__A2 (.I(_04523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09140__A2 (.I(_04523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09139__A2 (.I(_04523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09172__A2 (.I(_04533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09171__A2 (.I(_04533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09170__A2 (.I(_04533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09169__A2 (.I(_04533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09168__A2 (.I(_04533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09167__A2 (.I(_04533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09166__A2 (.I(_04533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09165__A2 (.I(_04533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09164__A2 (.I(_04533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09163__A2 (.I(_04533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09162__A2 (.I(_04533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09161__A2 (.I(_04533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09160__A2 (.I(_04533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09159__A2 (.I(_04533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09158__A2 (.I(_04533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09157__A2 (.I(_04533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09190__A2 (.I(_04543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09189__A2 (.I(_04543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09188__A2 (.I(_04543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09187__A2 (.I(_04543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09186__A2 (.I(_04543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09185__A2 (.I(_04543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09184__A2 (.I(_04543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09183__A2 (.I(_04543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09182__A2 (.I(_04543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09181__A2 (.I(_04543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09180__A2 (.I(_04543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09179__A2 (.I(_04543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09178__A2 (.I(_04543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09177__A2 (.I(_04543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09176__A2 (.I(_04543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09175__A2 (.I(_04543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09208__A2 (.I(_04553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09207__A2 (.I(_04553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09206__A2 (.I(_04553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09205__A2 (.I(_04553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09204__A2 (.I(_04553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09203__A2 (.I(_04553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09202__A2 (.I(_04553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09201__A2 (.I(_04553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09200__A2 (.I(_04553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09199__A2 (.I(_04553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09198__A2 (.I(_04553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09197__A2 (.I(_04553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09196__A2 (.I(_04553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09195__A2 (.I(_04553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09194__A2 (.I(_04553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09193__A2 (.I(_04553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09226__A2 (.I(_04563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09225__A2 (.I(_04563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09224__A2 (.I(_04563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09223__A2 (.I(_04563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09222__A2 (.I(_04563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09221__A2 (.I(_04563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09220__A2 (.I(_04563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09219__A2 (.I(_04563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09218__A2 (.I(_04563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09217__A2 (.I(_04563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09216__A2 (.I(_04563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09215__A2 (.I(_04563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09214__A2 (.I(_04563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09213__A2 (.I(_04563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09212__A2 (.I(_04563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09211__A2 (.I(_04563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09244__A2 (.I(_04573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09243__A2 (.I(_04573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09242__A2 (.I(_04573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09241__A2 (.I(_04573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09240__A2 (.I(_04573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09239__A2 (.I(_04573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09238__A2 (.I(_04573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09237__A2 (.I(_04573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09236__A2 (.I(_04573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09235__A2 (.I(_04573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09234__A2 (.I(_04573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09233__A2 (.I(_04573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09232__A2 (.I(_04573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09231__A2 (.I(_04573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09230__A2 (.I(_04573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09229__A2 (.I(_04573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09262__A2 (.I(_04583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09261__A2 (.I(_04583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09260__A2 (.I(_04583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09259__A2 (.I(_04583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09258__A2 (.I(_04583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09257__A2 (.I(_04583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09256__A2 (.I(_04583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09255__A2 (.I(_04583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09254__A2 (.I(_04583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09253__A2 (.I(_04583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09252__A2 (.I(_04583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09251__A2 (.I(_04583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09250__A2 (.I(_04583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09249__A2 (.I(_04583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09248__A2 (.I(_04583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09247__A2 (.I(_04583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09280__A2 (.I(_04593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09279__A2 (.I(_04593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09278__A2 (.I(_04593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09277__A2 (.I(_04593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09276__A2 (.I(_04593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09275__A2 (.I(_04593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09274__A2 (.I(_04593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09273__A2 (.I(_04593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09272__A2 (.I(_04593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09271__A2 (.I(_04593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09270__A2 (.I(_04593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09269__A2 (.I(_04593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09268__A2 (.I(_04593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09267__A2 (.I(_04593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09266__A2 (.I(_04593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09265__A2 (.I(_04593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09298__A2 (.I(_04603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09297__A2 (.I(_04603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09296__A2 (.I(_04603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09295__A2 (.I(_04603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09294__A2 (.I(_04603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09293__A2 (.I(_04603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09292__A2 (.I(_04603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09291__A2 (.I(_04603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09290__A2 (.I(_04603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09289__A2 (.I(_04603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09288__A2 (.I(_04603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09287__A2 (.I(_04603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09286__A2 (.I(_04603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09285__A2 (.I(_04603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09284__A2 (.I(_04603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09283__A2 (.I(_04603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09316__A2 (.I(_04613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09315__A2 (.I(_04613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09314__A2 (.I(_04613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09313__A2 (.I(_04613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09312__A2 (.I(_04613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09311__A2 (.I(_04613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09310__A2 (.I(_04613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09309__A2 (.I(_04613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09308__A2 (.I(_04613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09307__A2 (.I(_04613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09306__A2 (.I(_04613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09305__A2 (.I(_04613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09304__A2 (.I(_04613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09303__A2 (.I(_04613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09302__A2 (.I(_04613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09301__A2 (.I(_04613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09675__A1 (.I(_04622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09657__A1 (.I(_04622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09639__A1 (.I(_04622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09621__A1 (.I(_04622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09585__A1 (.I(_04622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09567__A1 (.I(_04622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09549__A1 (.I(_04622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09531__A1 (.I(_04622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09472__A1 (.I(_04622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09454__A1 (.I(_04622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09436__A1 (.I(_04622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09418__A1 (.I(_04622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09400__A1 (.I(_04622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09382__A1 (.I(_04622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09346__A1 (.I(_04622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09321__A1 (.I(_04622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09342__A2 (.I(_04624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09341__A2 (.I(_04624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09339__A2 (.I(_04624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09338__A2 (.I(_04624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09336__A2 (.I(_04624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09335__A2 (.I(_04624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09333__A2 (.I(_04624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09332__A2 (.I(_04624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09330__A2 (.I(_04624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09329__A2 (.I(_04624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09327__A2 (.I(_04624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09326__A2 (.I(_04624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09324__A2 (.I(_04624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09323__A2 (.I(_04624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09321__A2 (.I(_04624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09320__A2 (.I(_04624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09677__A1 (.I(_04626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09659__A1 (.I(_04626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09641__A1 (.I(_04626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09623__A1 (.I(_04626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09587__A1 (.I(_04626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09569__A1 (.I(_04626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09551__A1 (.I(_04626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09533__A1 (.I(_04626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09474__A1 (.I(_04626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09456__A1 (.I(_04626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09438__A1 (.I(_04626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09420__A1 (.I(_04626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09402__A1 (.I(_04626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09384__A1 (.I(_04626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09348__A1 (.I(_04626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09324__A1 (.I(_04626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09679__A1 (.I(_04628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09661__A1 (.I(_04628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09643__A1 (.I(_04628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09625__A1 (.I(_04628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09589__A1 (.I(_04628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09571__A1 (.I(_04628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09553__A1 (.I(_04628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09535__A1 (.I(_04628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09476__A1 (.I(_04628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09458__A1 (.I(_04628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09440__A1 (.I(_04628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09422__A1 (.I(_04628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09404__A1 (.I(_04628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09386__A1 (.I(_04628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09350__A1 (.I(_04628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09327__A1 (.I(_04628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09681__A1 (.I(_04630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09663__A1 (.I(_04630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09645__A1 (.I(_04630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09627__A1 (.I(_04630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09591__A1 (.I(_04630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09573__A1 (.I(_04630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09555__A1 (.I(_04630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09537__A1 (.I(_04630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09478__A1 (.I(_04630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09460__A1 (.I(_04630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09442__A1 (.I(_04630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09424__A1 (.I(_04630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09406__A1 (.I(_04630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09388__A1 (.I(_04630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09352__A1 (.I(_04630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09330__A1 (.I(_04630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09683__A1 (.I(_04632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09665__A1 (.I(_04632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09647__A1 (.I(_04632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09629__A1 (.I(_04632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09593__A1 (.I(_04632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09575__A1 (.I(_04632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09557__A1 (.I(_04632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09539__A1 (.I(_04632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09480__A1 (.I(_04632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09462__A1 (.I(_04632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09444__A1 (.I(_04632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09426__A1 (.I(_04632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09408__A1 (.I(_04632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09390__A1 (.I(_04632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09354__A1 (.I(_04632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09333__A1 (.I(_04632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09685__A1 (.I(_04634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09667__A1 (.I(_04634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09649__A1 (.I(_04634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09631__A1 (.I(_04634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09595__A1 (.I(_04634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09577__A1 (.I(_04634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09559__A1 (.I(_04634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09541__A1 (.I(_04634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09482__A1 (.I(_04634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09464__A1 (.I(_04634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09446__A1 (.I(_04634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09428__A1 (.I(_04634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09410__A1 (.I(_04634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09392__A1 (.I(_04634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09356__A1 (.I(_04634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09336__A1 (.I(_04634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09687__A1 (.I(_04636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09669__A1 (.I(_04636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09651__A1 (.I(_04636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09633__A1 (.I(_04636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09597__A1 (.I(_04636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09579__A1 (.I(_04636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09561__A1 (.I(_04636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09543__A1 (.I(_04636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09484__A1 (.I(_04636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09466__A1 (.I(_04636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09448__A1 (.I(_04636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09430__A1 (.I(_04636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09412__A1 (.I(_04636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09394__A1 (.I(_04636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09358__A1 (.I(_04636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09339__A1 (.I(_04636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09689__A1 (.I(_04638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09671__A1 (.I(_04638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09653__A1 (.I(_04638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09635__A1 (.I(_04638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09599__A1 (.I(_04638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09581__A1 (.I(_04638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09563__A1 (.I(_04638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09545__A1 (.I(_04638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09486__A1 (.I(_04638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09468__A1 (.I(_04638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09450__A1 (.I(_04638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09432__A1 (.I(_04638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09414__A1 (.I(_04638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09396__A1 (.I(_04638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09360__A1 (.I(_04638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09342__A1 (.I(_04638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09360__A2 (.I(_04641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09359__A2 (.I(_04641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09358__A2 (.I(_04641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09357__A2 (.I(_04641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09356__A2 (.I(_04641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09355__A2 (.I(_04641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09354__A2 (.I(_04641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09353__A2 (.I(_04641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09352__A2 (.I(_04641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09351__A2 (.I(_04641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09350__A2 (.I(_04641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09349__A2 (.I(_04641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09348__A2 (.I(_04641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09347__A2 (.I(_04641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09346__A2 (.I(_04641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09345__A2 (.I(_04641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09378__A2 (.I(_04651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09377__A2 (.I(_04651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09376__A2 (.I(_04651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09375__A2 (.I(_04651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09374__A2 (.I(_04651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09373__A2 (.I(_04651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09372__A2 (.I(_04651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09371__A2 (.I(_04651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09370__A2 (.I(_04651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09369__A2 (.I(_04651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09368__A2 (.I(_04651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09367__A2 (.I(_04651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09366__A2 (.I(_04651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09365__A2 (.I(_04651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09364__A2 (.I(_04651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09363__A2 (.I(_04651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09380__I (.I(_04660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09396__A2 (.I(_04661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09395__A2 (.I(_04661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09394__A2 (.I(_04661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09393__A2 (.I(_04661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09392__A2 (.I(_04661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09391__A2 (.I(_04661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09390__A2 (.I(_04661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09389__A2 (.I(_04661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09388__A2 (.I(_04661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09387__A2 (.I(_04661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09386__A2 (.I(_04661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09385__A2 (.I(_04661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09384__A2 (.I(_04661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09383__A2 (.I(_04661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09382__A2 (.I(_04661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09381__A2 (.I(_04661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09414__A2 (.I(_04671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09413__A2 (.I(_04671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09412__A2 (.I(_04671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09411__A2 (.I(_04671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09410__A2 (.I(_04671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09409__A2 (.I(_04671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09408__A2 (.I(_04671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09407__A2 (.I(_04671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09406__A2 (.I(_04671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09405__A2 (.I(_04671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09404__A2 (.I(_04671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09403__A2 (.I(_04671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09402__A2 (.I(_04671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09401__A2 (.I(_04671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09400__A2 (.I(_04671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09399__A2 (.I(_04671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09416__I (.I(_04680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09432__A2 (.I(_04681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09431__A2 (.I(_04681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09430__A2 (.I(_04681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09429__A2 (.I(_04681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09428__A2 (.I(_04681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09427__A2 (.I(_04681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09426__A2 (.I(_04681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09425__A2 (.I(_04681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09424__A2 (.I(_04681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09423__A2 (.I(_04681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09422__A2 (.I(_04681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09421__A2 (.I(_04681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09420__A2 (.I(_04681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09419__A2 (.I(_04681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09418__A2 (.I(_04681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09417__A2 (.I(_04681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09450__A2 (.I(_04691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09449__A2 (.I(_04691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09448__A2 (.I(_04691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09447__A2 (.I(_04691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09446__A2 (.I(_04691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09445__A2 (.I(_04691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09444__A2 (.I(_04691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09443__A2 (.I(_04691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09442__A2 (.I(_04691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09441__A2 (.I(_04691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09440__A2 (.I(_04691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09439__A2 (.I(_04691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09438__A2 (.I(_04691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09437__A2 (.I(_04691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09436__A2 (.I(_04691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09435__A2 (.I(_04691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09468__A2 (.I(_04701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09467__A2 (.I(_04701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09466__A2 (.I(_04701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09465__A2 (.I(_04701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09464__A2 (.I(_04701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09463__A2 (.I(_04701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09462__A2 (.I(_04701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09461__A2 (.I(_04701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09460__A2 (.I(_04701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09459__A2 (.I(_04701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09458__A2 (.I(_04701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09457__A2 (.I(_04701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09456__A2 (.I(_04701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09455__A2 (.I(_04701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09454__A2 (.I(_04701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09453__A2 (.I(_04701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09486__A2 (.I(_04711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09485__A2 (.I(_04711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09484__A2 (.I(_04711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09483__A2 (.I(_04711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09482__A2 (.I(_04711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09481__A2 (.I(_04711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09480__A2 (.I(_04711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09479__A2 (.I(_04711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09478__A2 (.I(_04711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09477__A2 (.I(_04711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09476__A2 (.I(_04711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09475__A2 (.I(_04711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09474__A2 (.I(_04711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09473__A2 (.I(_04711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09472__A2 (.I(_04711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09471__A2 (.I(_04711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09506__A2 (.I(_04723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09505__B (.I(_04723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09503__S (.I(_04723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09500__A2 (.I(_04723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09499__A1 (.I(_04723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09496__A2 (.I(_04723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09495__A1 (.I(_04723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09545__A2 (.I(_04752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09544__A2 (.I(_04752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09543__A2 (.I(_04752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09542__A2 (.I(_04752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09541__A2 (.I(_04752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09540__A2 (.I(_04752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09539__A2 (.I(_04752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09538__A2 (.I(_04752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09537__A2 (.I(_04752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09536__A2 (.I(_04752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09535__A2 (.I(_04752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09534__A2 (.I(_04752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09533__A2 (.I(_04752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09532__A2 (.I(_04752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09531__A2 (.I(_04752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09530__A2 (.I(_04752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09563__A2 (.I(_04762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09562__A2 (.I(_04762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09561__A2 (.I(_04762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09560__A2 (.I(_04762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09559__A2 (.I(_04762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09558__A2 (.I(_04762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09557__A2 (.I(_04762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09556__A2 (.I(_04762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09555__A2 (.I(_04762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09554__A2 (.I(_04762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09553__A2 (.I(_04762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09552__A2 (.I(_04762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09551__A2 (.I(_04762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09550__A2 (.I(_04762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09549__A2 (.I(_04762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09548__A2 (.I(_04762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09581__A2 (.I(_04772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09580__A2 (.I(_04772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09579__A2 (.I(_04772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09578__A2 (.I(_04772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09577__A2 (.I(_04772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09576__A2 (.I(_04772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09575__A2 (.I(_04772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09574__A2 (.I(_04772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09573__A2 (.I(_04772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09572__A2 (.I(_04772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09571__A2 (.I(_04772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09570__A2 (.I(_04772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09569__A2 (.I(_04772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09568__A2 (.I(_04772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09567__A2 (.I(_04772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09566__A2 (.I(_04772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09599__A2 (.I(_04782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09598__A2 (.I(_04782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09597__A2 (.I(_04782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09596__A2 (.I(_04782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09595__A2 (.I(_04782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09594__A2 (.I(_04782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09593__A2 (.I(_04782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09592__A2 (.I(_04782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09591__A2 (.I(_04782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09590__A2 (.I(_04782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09589__A2 (.I(_04782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09588__A2 (.I(_04782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09587__A2 (.I(_04782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09586__A2 (.I(_04782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09585__A2 (.I(_04782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09584__A2 (.I(_04782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09617__A2 (.I(_04792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09616__A2 (.I(_04792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09615__A2 (.I(_04792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09614__A2 (.I(_04792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09613__A2 (.I(_04792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09612__A2 (.I(_04792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09611__A2 (.I(_04792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09610__A2 (.I(_04792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09609__A2 (.I(_04792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09608__A2 (.I(_04792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09607__A2 (.I(_04792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09606__A2 (.I(_04792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09605__A2 (.I(_04792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09604__A2 (.I(_04792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09603__A2 (.I(_04792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09602__A2 (.I(_04792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09635__A2 (.I(_04802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09634__A2 (.I(_04802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09633__A2 (.I(_04802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09632__A2 (.I(_04802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09631__A2 (.I(_04802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09630__A2 (.I(_04802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09629__A2 (.I(_04802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09628__A2 (.I(_04802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09627__A2 (.I(_04802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09626__A2 (.I(_04802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09625__A2 (.I(_04802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09624__A2 (.I(_04802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09623__A2 (.I(_04802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09622__A2 (.I(_04802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09621__A2 (.I(_04802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09620__A2 (.I(_04802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09653__A2 (.I(_04812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09652__A2 (.I(_04812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09651__A2 (.I(_04812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09650__A2 (.I(_04812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09649__A2 (.I(_04812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09648__A2 (.I(_04812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09647__A2 (.I(_04812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09646__A2 (.I(_04812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09645__A2 (.I(_04812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09644__A2 (.I(_04812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09643__A2 (.I(_04812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09642__A2 (.I(_04812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09641__A2 (.I(_04812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09640__A2 (.I(_04812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09639__A2 (.I(_04812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09638__A2 (.I(_04812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09671__A2 (.I(_04822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09670__A2 (.I(_04822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09669__A2 (.I(_04822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09668__A2 (.I(_04822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09667__A2 (.I(_04822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09666__A2 (.I(_04822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09665__A2 (.I(_04822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09664__A2 (.I(_04822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09663__A2 (.I(_04822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09662__A2 (.I(_04822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09661__A2 (.I(_04822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09660__A2 (.I(_04822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09659__A2 (.I(_04822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09658__A2 (.I(_04822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09657__A2 (.I(_04822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09656__A2 (.I(_04822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09689__A2 (.I(_04832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09688__A2 (.I(_04832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09687__A2 (.I(_04832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09686__A2 (.I(_04832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09685__A2 (.I(_04832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09684__A2 (.I(_04832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09683__A2 (.I(_04832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09682__A2 (.I(_04832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09681__A2 (.I(_04832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09680__A2 (.I(_04832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09679__A2 (.I(_04832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09678__A2 (.I(_04832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09677__A2 (.I(_04832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09676__A2 (.I(_04832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09675__A2 (.I(_04832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09674__A2 (.I(_04832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11114__CLK (.I(io_in[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11113__CLK (.I(io_in[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11112__CLK (.I(io_in[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11111__CLK (.I(io_in[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11110__CLK (.I(io_in[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11109__CLK (.I(io_in[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11108__CLK (.I(io_in[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11107__CLK (.I(io_in[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11106__CLK (.I(io_in[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11104__CLK (.I(io_in[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11105__CLK (.I(io_in[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11093__CLK (.I(io_in[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11094__CLK (.I(io_in[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11103__CLK (.I(io_in[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11095__CLK (.I(io_in[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11102__CLK (.I(io_in[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11101__CLK (.I(io_in[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11100__CLK (.I(io_in[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11119__CLK (.I(io_in[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11099__CLK (.I(io_in[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11098__CLK (.I(io_in[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11097__CLK (.I(io_in[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11096__CLK (.I(io_in[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11118__CLK (.I(io_in[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11117__CLK (.I(io_in[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11116__CLK (.I(io_in[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11115__CLK (.I(io_in[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11089__CLK (.I(io_in[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11088__CLK (.I(io_in[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11092__CLK (.I(io_in[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11091__CLK (.I(io_in[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11120__CLK (.I(io_in[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11121__CLK (.I(io_in[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11122__CLK (.I(io_in[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11125__CLK (.I(io_in[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11124__CLK (.I(io_in[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11127__CLK (.I(io_in[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11126__CLK (.I(io_in[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11090__CLK (.I(io_in[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11123__CLK (.I(io_in[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11132__CLK (.I(io_in[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11131__CLK (.I(io_in[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11130__CLK (.I(io_in[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11145__CLK (.I(io_in[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11137__CLK (.I(io_in[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11140__CLK (.I(io_in[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11141__CLK (.I(io_in[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11143__CLK (.I(io_in[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11136__CLK (.I(io_in[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11135__CLK (.I(io_in[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11142__CLK (.I(io_in[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11138__CLK (.I(io_in[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11139__CLK (.I(io_in[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11144__CLK (.I(io_in[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11134__CLK (.I(io_in[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11133__CLK (.I(io_in[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11153__CLK (.I(io_in[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11154__CLK (.I(io_in[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11152__CLK (.I(io_in[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11149__CLK (.I(io_in[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11148__CLK (.I(io_in[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11087__CLKN (.I(io_in[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11166__I (.I(io_in[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11157__CLK (.I(io_in[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11151__CLK (.I(io_in[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11150__CLK (.I(io_in[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11147__CLK (.I(io_in[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11146__CLK (.I(io_in[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11129__CLK (.I(io_in[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11128__CLK (.I(io_in[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11155__CLK (.I(io_in[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11156__CLK (.I(io_in[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05835__I (.I(io_in[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05830__A1 (.I(io_in[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05828__I (.I(io_in[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10497__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10928__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10925__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10494__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10207__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10206__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10119__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10303__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10159__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10498__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10929__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10118__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10302__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10158__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10111__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10489__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10924__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10493__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10490__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10205__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10117__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10301__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10157__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10107__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10486__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10112__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10108__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10487__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10110__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10496__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10927__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10109__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10495__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10488__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10926__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09954__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09757__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10155__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10299__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10044__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09948__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09751__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09952__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09755__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10048__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09859__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10115__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10203__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10485__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10043__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09756__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09953__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10249__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10233__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10217__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09860__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09861__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10050__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10049__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09855__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09857__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09951__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09950__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09753__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09754__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10046__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09856__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09752__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09858__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10045__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10047__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09949__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09854__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09947__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09750__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10734__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11026__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10737__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10736__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10729__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10728__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09745__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09746__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10208__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10120__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10304__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10160__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10209__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10121__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10161__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10305__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10725__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10156__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10300__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10735__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10727__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10733__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10726__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10210__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09743__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11024__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09744__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10204__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10116__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10173__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10165__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10738__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10730__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09747__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10739__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09941__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11025__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09927__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10163__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10174__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09943__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10166__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09923__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10171__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09942__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09925__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09939__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10172__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09940__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09924__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10167__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09928__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11023__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11027__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10175__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11028__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09748__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10731__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10500__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10931__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10492__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10114__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09742__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10306__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11022__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10162__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10122__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10491__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10113__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10499__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10930__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10227__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09911__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10211__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10213__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10229__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10245__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09907__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09909__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10216__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10248__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10232__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10231__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10247__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10215__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10192__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09945__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09929__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09930__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10176__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10168__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11029__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09749__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10164__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09944__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10732__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10740__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10293__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10186__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10298__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10194__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09912__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09914__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09946__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10178__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10177__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10170__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10169__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09913__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10277__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10264__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10256__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10271__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10263__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10255__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10244__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10243__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10212__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10280__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10272__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10269__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10261__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10253__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10196__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10153__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10138__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10266__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10262__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10258__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10274__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10254__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10201__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10137__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10202__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10146__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10282__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10270__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10145__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10279__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10557__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10555__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10554__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10556__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10268__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10267__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10275__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10257__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10252__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10265__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10260__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10259__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10251__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10276__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10281__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10273__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10560__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10796__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10810__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10801__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10799__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10559__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10558__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10800__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10809__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10802__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10553__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10552__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10551__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10154__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10278__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10197__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10195__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10133__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10797__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10149__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10798__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10141__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10621__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10620__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10214__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09910__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10230__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10246__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10289__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10297__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10234__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10250__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09908__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10218__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10228__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09900__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10150__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10142__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10148__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10140__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09905__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10321__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10296__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10295__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09901__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09903__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10287__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10285__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10322__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10317__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09906__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10290__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10291__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10318__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10294__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09899__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10288__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10315__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10320__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09707__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10283__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09904__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09708__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09704__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10286__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09902__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10134__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10198__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10132__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10292__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10284__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10129__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10124__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10360__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10144__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10143__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10123__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11072__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10130__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10136__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10200__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10135__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10199__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10131__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10139__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10363__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10356__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10367__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11073__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10152__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11075__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10362__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10355__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10151__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10619__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10618__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10361__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11071__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10147__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09759__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10316__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09706__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09703__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09702__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09709__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09719__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11054__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10127__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10128__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10126__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10125__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10359__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11080__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11081__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10364__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10365__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10358__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10357__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11068__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11067__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11066__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11069__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10366__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10182__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10189__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10190__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09983__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10181__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09975__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09967__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09991__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09926__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09972__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09964__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09976__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09984__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09968__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09992__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09988__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10187__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09980__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10904__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09959__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10183__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10191__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10902__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10903__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09955__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10900__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09958__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09957__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09726__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09877__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10179__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09971__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09969__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09963__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09973__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09965__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09989__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09981__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09978__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09970__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09994__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09919__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09977__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09985__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09993__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09986__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09974__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09966__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09916__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09982__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09990__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10853__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09767__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09728__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09730__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10856__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09770__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09935__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09979__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09987__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10184__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10905__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09960__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10901__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09733__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09732__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09727__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10035__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09867__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09956__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09875__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09869__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09961__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10185__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10193__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09868__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10859__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09922__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09773__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09938__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09871__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09879__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09878__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09729__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10038__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10039__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09932__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09715__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09739__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09740__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09741__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09731__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09876__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09873__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10906__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09874__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09881__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09882__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11062__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11061__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09717__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09716__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09872__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09870__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09880__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09936__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09920__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09772__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11004__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10996__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11021__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11013__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09921__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11020__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11012__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11005__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10997__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10858__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09937__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09712__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09736__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10999__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10991__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11007__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11015__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11010__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09738__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11057__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11060__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11059__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09714__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11006__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11014__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11016__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11000__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10998__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10990__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10992__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11008__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10995__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11009__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11017__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10993__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11001__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11019__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11011__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11003__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09771__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09766__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10857__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10855__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10852__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09931__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09934__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09918__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09769__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09915__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09933__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10854__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09917__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09768__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10994__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11018__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10188__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10180__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11002__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09997__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10002__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10042__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10041__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10037__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10680__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10638__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10681__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10639__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10001__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09962__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10907__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10036__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10319__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09760__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09761__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09724__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09723__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10795__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10794__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10632__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10674__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09995__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10886__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10887__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09721__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09720__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10890__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10889__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09705__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10676__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10634__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10679__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09735__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09734__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09710__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10314__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10313__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10040__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11056__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11055__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09711__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10770__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10312__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10790__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10793__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10307__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10637__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10000__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10308__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10636__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10678__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09718__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09725__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09722__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09764__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10884__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10885__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09996__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09763__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10891__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10633__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10789__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10888__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10788__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09828__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09780__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09820__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09818__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09758__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09762__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09765__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09827__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09779__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09826__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09778__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10741__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09998__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10422__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10635__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10791__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10414__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10418__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10675__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10677__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10792__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09999__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09814__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11052__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10978__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10979__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11053__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10419__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10411__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10974__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11048__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09822__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09774__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10423__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10415__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10410__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10435__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10765__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10309__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10747__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10743__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10776__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10772__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10431__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10768__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10764__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10311__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09737__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09713__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11058__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10746__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10762__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10775__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10310__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10434__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10769__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10744__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10773__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10766__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10763__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10432__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10771__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10767__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10938__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10934__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10914__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10948__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10964__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10932__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10908__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10971__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10915__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10939__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10954__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10970__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10966__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10955__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10950__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10965__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10967__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10937__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10936__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10935__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10933__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10911__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10910__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10949__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10969__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10968__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10952__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10953__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10951__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10722__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10898__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10429__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10777__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10947__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10742__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10436__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10430__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10748__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10420__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10745__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10774__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10433__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10719__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10956__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10723__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10940__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10899__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11050__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10716__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10892__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10874__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10976__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10963__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10412__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10897__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10720__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10721__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10962__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10960__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10944__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10945__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10946__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10961__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10896__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10913__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10912__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10909__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10893__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10943__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10958__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10942__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10869__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10870__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10894__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10957__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10941__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10872__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10717__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10895__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10718__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10959__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10549__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10808__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10806__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10804__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10803__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10807__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10562__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10561__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10550__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10610__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10609__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10805__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10564__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10563__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10988__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10607__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10613__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10612__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10583__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10615__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10608__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10585__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10614__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10606__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10616__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10750__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10605__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10617__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10542__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10611__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10567__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10811__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10547__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10546__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10565__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10566__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10568__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10569__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10548__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10543__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10545__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10544__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10400__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10671__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10426__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10622__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10581__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10724__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10584__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10786__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10588__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10582__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10587__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10586__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10640__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10603__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11084__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10752__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10751__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09864__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09865__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09866__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11076__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09863__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10749__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10753__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10604__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10602__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10600__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09848__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11085__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10238__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10377__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10220__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11079__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11065__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11064__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11077__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11078__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10236__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11082__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11083__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11070__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10386__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10237__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10393__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10382__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10225__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10240__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10241__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09852__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09849__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10378__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10385__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10221__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09846__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10590__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10589__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09808__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09832__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10982__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10983__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10981__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09806__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10235__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10239__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10986__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10623__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10984__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10980__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09850__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10383__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10226__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10381__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10224__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09812__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09836__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09853__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09813__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09833__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09809__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10398__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10390__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10242__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09835__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09811__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09837__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09830__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10987__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10985__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10425__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09810__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10389__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09851__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09807__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09847__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10397__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10399__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10058__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10601__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10591__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11086__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10691__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10688__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10689__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10570__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10687__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10686__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10787__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10685__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10571__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10572__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10541__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10645__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10644__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10643__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10690__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10713__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10712__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10424__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10428__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11063__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10682__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10683__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10641__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10672__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10673__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10684__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10670__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10714__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10715__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10642__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10648__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10699__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10696__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10697__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10646__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10693__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10692__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10695__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10694__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10647__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10698__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10654__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10656__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10650__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10651__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10652__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10711__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10706__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10705__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10708__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10707__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10703__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10704__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10700__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10701__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10702__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10710__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10709__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10663__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10661__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10660__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10658__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10655__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10649__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10653__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10662__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10659__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10657__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10004__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10012__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10401__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10402__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10403__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10021__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10005__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10989__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10407__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10013__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10406__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10427__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09834__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10668__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10028__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10014__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10006__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10020__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10011__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09862__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10405__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10019__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11074__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10404__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10027__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10003__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10015__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10669__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10029__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10084__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10051__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10074__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10077__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10085__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10101__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10093__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09831__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10066__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10443__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10087__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10078__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10059__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10099__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10091__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10083__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10092__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10100__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10086__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10067__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10076__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10075__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10666__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10665__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10030__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10008__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10016__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10667__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10031__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10023__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10010__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10009__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10018__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10017__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10022__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10007__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10664__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10032__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10438__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10082__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10081__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10079__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10089__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10090__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10103__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10095__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10094__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10088__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10080__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10102__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10098__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10106__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10105__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10097__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10033__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10034__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10025__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10026__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10024__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10096__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10104__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09823__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09775__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09781__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09829__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09776__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09824__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10222__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10379__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09889__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09888__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09819__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09887__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09788__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09844__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09796__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10376__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09789__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09885__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09816__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10395__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10394__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09821__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09815__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09890__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09884__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10387__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09817__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09886__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10409__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11047__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10416__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09883__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09825__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09777__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11046__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10408__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11049__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10417__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10975__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09897__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09894__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09893__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09785__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09784__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09840__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09841__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09801__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09793__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09792__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10973__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10972__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09787__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09804__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10392__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10384__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10380__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10223__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09797__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09805__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09845__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10219__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10391__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10056__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10057__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10922__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10923__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10396__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09786__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10460__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09898__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09891__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09838__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09782__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09798__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09790__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10476__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10469__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10453__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10525__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09800__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09839__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09791__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09799__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09783__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10474__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09896__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09895__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10471__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09892__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09842__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09794__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09802__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10532__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10388__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09843__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09795__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09803__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10918__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10921__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10876__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10882__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11051__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10860__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10843__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10836__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10867__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10866__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10842__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10421__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10413__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10868__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10883__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10875__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10834__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10818__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10827__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10835__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10831__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10826__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10819__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10828__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10820__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10977__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10863__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10877__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10840__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10861__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10878__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10865__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10864__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10862__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10837__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10839__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10841__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10880__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10879__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10871__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10881__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10873__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10830__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10838__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10817__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10816__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10833__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10832__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10824__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10825__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10822__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10829__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10821__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10823__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10531__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10851__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11037__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10844__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10785__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11030__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10475__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10459__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10784__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10850__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11044__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10812__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10815__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11038__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11045__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10757__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10754__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10472__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10374__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10375__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10516__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10456__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10528__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10473__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10515__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10778__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10761__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10760__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11042__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11031__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10845__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10779__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10846__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11032__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10780__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11036__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11043__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11040__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10814__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10813__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11039__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11041__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11034__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10849__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11035__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10783__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10781__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10848__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10782__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10755__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10847__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11033__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10756__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10919__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10072__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10073__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10065__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10920__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10917__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10916__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10053__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10063__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10062__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10055__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10054__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10052__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10064__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10445__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10070__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10071__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10069__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10068__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10060__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10447__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10439__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10451__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10437__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10539__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10061__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10458__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10530__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10455__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10454__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10527__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10526__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10470__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10592__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10333__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10337__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10329__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10353__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10327__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10335__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10325__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10345__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10535__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10626__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10534__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10625__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10444__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10452__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10446__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10442__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10449__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10441__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10440__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10448__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10450__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10533__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10624__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10630__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10537__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10628__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10629__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10631__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10627__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10536__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10540__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10538__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10593__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10502__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10599__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10501__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10338__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10346__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10330__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10351__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10334__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10323__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10354__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10347__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10339__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10331__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10508__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10340__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10342__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10348__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10350__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10344__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10352__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10326__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10336__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10324__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10328__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10332__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10349__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10341__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10343__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10373__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10463__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10468__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10509__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10457__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10512__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10372__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10371__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10370__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10369__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10368__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10529__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10510__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10484__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10467__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10483__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10477__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10461__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10480__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10464__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10598__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10594__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10519__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10517__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10579__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10523__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10462__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10478__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10482__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10481__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10479__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10513__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10514__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10466__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10465__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10759__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10758__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10511__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10521__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10522__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10503__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10575__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10595__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10597__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10596__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10507__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10574__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10520__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10504__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10576__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10518__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10573__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10577__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10578__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10505__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10506__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10524__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10580__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08714__I0 (.I(\u_arbiter.i_wb_cpu_dbus_adr[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08712__I1 (.I(\u_arbiter.i_wb_cpu_dbus_adr[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06003__B2 (.I(\u_arbiter.i_wb_cpu_dbus_adr[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08758__A1 (.I(\u_arbiter.i_wb_cpu_dbus_adr[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08690__I0 (.I(\u_arbiter.i_wb_cpu_dbus_adr[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05949__C2 (.I(\u_arbiter.i_wb_cpu_dbus_adr[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08752__I0 (.I(\u_arbiter.i_wb_cpu_dbus_adr[31] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08750__A2 (.I(\u_arbiter.i_wb_cpu_dbus_adr[31] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08746__I1 (.I(\u_arbiter.i_wb_cpu_dbus_adr[31] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06092__B2 (.I(\u_arbiter.i_wb_cpu_dbus_adr[31] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08696__I0 (.I(\u_arbiter.i_wb_cpu_dbus_adr[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08694__I1 (.I(\u_arbiter.i_wb_cpu_dbus_adr[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05962__B2 (.I(\u_arbiter.i_wb_cpu_dbus_adr[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08700__I0 (.I(\u_arbiter.i_wb_cpu_dbus_adr[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08698__I1 (.I(\u_arbiter.i_wb_cpu_dbus_adr[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05970__B2 (.I(\u_arbiter.i_wb_cpu_dbus_adr[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08151__A2 (.I(\u_arbiter.i_wb_cpu_dbus_dat[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08144__A1 (.I(\u_arbiter.i_wb_cpu_dbus_dat[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08141__B2 (.I(\u_arbiter.i_wb_cpu_dbus_dat[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08135__A1 (.I(\u_arbiter.i_wb_cpu_dbus_dat[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06592__A3 (.I(\u_arbiter.i_wb_cpu_dbus_dat[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05863__A1 (.I(\u_arbiter.i_wb_cpu_dbus_dat[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05781__I0 (.I(\u_arbiter.i_wb_cpu_dbus_dat[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08186__A1 (.I(\u_arbiter.i_wb_cpu_dbus_dat[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08184__B2 (.I(\u_arbiter.i_wb_cpu_dbus_dat[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05884__I1 (.I(\u_arbiter.i_wb_cpu_dbus_dat[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08204__A1 (.I(\u_arbiter.i_wb_cpu_dbus_dat[16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08202__B2 (.I(\u_arbiter.i_wb_cpu_dbus_dat[16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05897__I1 (.I(\u_arbiter.i_wb_cpu_dbus_dat[16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05781__I2 (.I(\u_arbiter.i_wb_cpu_dbus_dat[16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08213__A1 (.I(\u_arbiter.i_wb_cpu_dbus_dat[19] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08211__B2 (.I(\u_arbiter.i_wb_cpu_dbus_dat[19] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05903__I1 (.I(\u_arbiter.i_wb_cpu_dbus_dat[19] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08151__A3 (.I(\u_arbiter.i_wb_cpu_dbus_dat[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08146__A1 (.I(\u_arbiter.i_wb_cpu_dbus_dat[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08144__A2 (.I(\u_arbiter.i_wb_cpu_dbus_dat[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08137__A1 (.I(\u_arbiter.i_wb_cpu_dbus_dat[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06592__A4 (.I(\u_arbiter.i_wb_cpu_dbus_dat[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05866__I1 (.I(\u_arbiter.i_wb_cpu_dbus_dat[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08219__A1 (.I(\u_arbiter.i_wb_cpu_dbus_dat[21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08217__B2 (.I(\u_arbiter.i_wb_cpu_dbus_dat[21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05907__I1 (.I(\u_arbiter.i_wb_cpu_dbus_dat[21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08229__B2 (.I(\u_arbiter.i_wb_cpu_dbus_dat[24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08226__B2 (.I(\u_arbiter.i_wb_cpu_dbus_dat[24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05913__I1 (.I(\u_arbiter.i_wb_cpu_dbus_dat[24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05781__I3 (.I(\u_arbiter.i_wb_cpu_dbus_dat[24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08239__A1 (.I(\u_arbiter.i_wb_cpu_dbus_dat[28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08237__B2 (.I(\u_arbiter.i_wb_cpu_dbus_dat[28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05922__I1 (.I(\u_arbiter.i_wb_cpu_dbus_dat[28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08153__A1 (.I(\u_arbiter.i_wb_cpu_dbus_dat[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08151__A1 (.I(\u_arbiter.i_wb_cpu_dbus_dat[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08143__A1 (.I(\u_arbiter.i_wb_cpu_dbus_dat[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06592__A2 (.I(\u_arbiter.i_wb_cpu_dbus_dat[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05868__I1 (.I(\u_arbiter.i_wb_cpu_dbus_dat[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08167__B2 (.I(\u_arbiter.i_wb_cpu_dbus_dat[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08162__A1 (.I(\u_arbiter.i_wb_cpu_dbus_dat[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08158__A1 (.I(\u_arbiter.i_wb_cpu_dbus_dat[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06593__A1 (.I(\u_arbiter.i_wb_cpu_dbus_dat[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05872__I1 (.I(\u_arbiter.i_wb_cpu_dbus_dat[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08171__A1 (.I(\u_arbiter.i_wb_cpu_dbus_dat[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08166__A1 (.I(\u_arbiter.i_wb_cpu_dbus_dat[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06594__A1 (.I(\u_arbiter.i_wb_cpu_dbus_dat[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05874__I1 (.I(\u_arbiter.i_wb_cpu_dbus_dat[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05740__A2 (.I(\u_arbiter.i_wb_cpu_dbus_dat[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08174__A1 (.I(\u_arbiter.i_wb_cpu_dbus_dat[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06597__A1 (.I(\u_arbiter.i_wb_cpu_dbus_dat[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05876__I1 (.I(\u_arbiter.i_wb_cpu_dbus_dat[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08180__A1 (.I(\u_arbiter.i_wb_cpu_dbus_dat[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08178__B2 (.I(\u_arbiter.i_wb_cpu_dbus_dat[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05880__I1 (.I(\u_arbiter.i_wb_cpu_dbus_dat[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05781__I1 (.I(\u_arbiter.i_wb_cpu_dbus_dat[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08497__A3 (.I(\u_arbiter.i_wb_cpu_dbus_we ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06118__A2 (.I(\u_arbiter.i_wb_cpu_dbus_we ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05841__I (.I(\u_arbiter.i_wb_cpu_dbus_we ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05751__A2 (.I(\u_arbiter.i_wb_cpu_dbus_we ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05700__S (.I(\u_arbiter.i_wb_cpu_dbus_we ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05691__A1 (.I(\u_arbiter.i_wb_cpu_dbus_we ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05690__A1 (.I(\u_arbiter.i_wb_cpu_dbus_we ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05684__A1 (.I(\u_arbiter.i_wb_cpu_dbus_we ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08784__A1 (.I(\u_arbiter.i_wb_cpu_ibus_adr[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06112__A2 (.I(\u_arbiter.i_wb_cpu_ibus_adr[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05935__A1 (.I(\u_arbiter.i_wb_cpu_ibus_adr[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05788__A2 (.I(\u_arbiter.i_wb_cpu_ibus_adr[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05755__B (.I(\u_arbiter.i_wb_cpu_ibus_adr[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05728__A1 (.I(\u_arbiter.i_wb_cpu_ibus_adr[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09047__A1 (.I(\u_arbiter.i_wb_cpu_ibus_adr[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08786__A1 (.I(\u_arbiter.i_wb_cpu_ibus_adr[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08784__B2 (.I(\u_arbiter.i_wb_cpu_ibus_adr[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08266__A2 (.I(\u_arbiter.i_wb_cpu_ibus_adr[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06586__A2 (.I(\u_arbiter.i_wb_cpu_ibus_adr[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05938__A1 (.I(\u_arbiter.i_wb_cpu_ibus_adr[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08594__I1 (.I(\u_arbiter.i_wb_cpu_rdt[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08286__A2 (.I(\u_arbiter.i_wb_cpu_rdt[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08272__I0 (.I(\u_arbiter.i_wb_cpu_rdt[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08141__A1 (.I(\u_arbiter.i_wb_cpu_rdt[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05853__A1 (.I(\u_arbiter.i_wb_cpu_rdt[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08441__I1 (.I(\u_arbiter.i_wb_cpu_rdt[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08374__A2 (.I(\u_arbiter.i_wb_cpu_rdt[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08295__I0 (.I(\u_arbiter.i_wb_cpu_rdt[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08187__A1 (.I(\u_arbiter.i_wb_cpu_rdt[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05878__I0 (.I(\u_arbiter.i_wb_cpu_rdt[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08512__I1 (.I(\u_arbiter.i_wb_cpu_rdt[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08293__A2 (.I(\u_arbiter.i_wb_cpu_rdt[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08190__A1 (.I(\u_arbiter.i_wb_cpu_rdt[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05880__I0 (.I(\u_arbiter.i_wb_cpu_rdt[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08525__I1 (.I(\u_arbiter.i_wb_cpu_rdt[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08378__I0 (.I(\u_arbiter.i_wb_cpu_rdt[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08307__A2 (.I(\u_arbiter.i_wb_cpu_rdt[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08193__A1 (.I(\u_arbiter.i_wb_cpu_rdt[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05882__I0 (.I(\u_arbiter.i_wb_cpu_rdt[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08532__I1 (.I(\u_arbiter.i_wb_cpu_rdt[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08347__I0 (.I(\u_arbiter.i_wb_cpu_rdt[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08289__A2 (.I(\u_arbiter.i_wb_cpu_rdt[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08196__A1 (.I(\u_arbiter.i_wb_cpu_rdt[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05884__I0 (.I(\u_arbiter.i_wb_cpu_rdt[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08538__I1 (.I(\u_arbiter.i_wb_cpu_rdt[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08349__A2 (.I(\u_arbiter.i_wb_cpu_rdt[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08277__I0 (.I(\u_arbiter.i_wb_cpu_rdt[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08199__A1 (.I(\u_arbiter.i_wb_cpu_rdt[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05886__I0 (.I(\u_arbiter.i_wb_cpu_rdt[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08643__I1 (.I(\u_arbiter.i_wb_cpu_rdt[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08319__I0 (.I(\u_arbiter.i_wb_cpu_rdt[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08280__A2 (.I(\u_arbiter.i_wb_cpu_rdt[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08202__A1 (.I(\u_arbiter.i_wb_cpu_rdt[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05888__I0 (.I(\u_arbiter.i_wb_cpu_rdt[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09069__I0 (.I(\u_arbiter.i_wb_cpu_rdt[16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08594__I0 (.I(\u_arbiter.i_wb_cpu_rdt[16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08205__A1 (.I(\u_arbiter.i_wb_cpu_rdt[16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05891__I0 (.I(\u_arbiter.i_wb_cpu_rdt[16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09071__I0 (.I(\u_arbiter.i_wb_cpu_rdt[17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08611__A2 (.I(\u_arbiter.i_wb_cpu_rdt[17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08208__A1 (.I(\u_arbiter.i_wb_cpu_rdt[17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05893__I0 (.I(\u_arbiter.i_wb_cpu_rdt[17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09073__I0 (.I(\u_arbiter.i_wb_cpu_rdt[18] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08627__A2 (.I(\u_arbiter.i_wb_cpu_rdt[18] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08211__A1 (.I(\u_arbiter.i_wb_cpu_rdt[18] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05895__I0 (.I(\u_arbiter.i_wb_cpu_rdt[18] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09075__I0 (.I(\u_arbiter.i_wb_cpu_rdt[19] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08636__A2 (.I(\u_arbiter.i_wb_cpu_rdt[19] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08214__A1 (.I(\u_arbiter.i_wb_cpu_rdt[19] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05897__I0 (.I(\u_arbiter.i_wb_cpu_rdt[19] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09077__I0 (.I(\u_arbiter.i_wb_cpu_rdt[20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08390__I0 (.I(\u_arbiter.i_wb_cpu_rdt[20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08217__A1 (.I(\u_arbiter.i_wb_cpu_rdt[20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05899__I0 (.I(\u_arbiter.i_wb_cpu_rdt[20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09079__I0 (.I(\u_arbiter.i_wb_cpu_rdt[21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08401__I0 (.I(\u_arbiter.i_wb_cpu_rdt[21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08220__A1 (.I(\u_arbiter.i_wb_cpu_rdt[21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05901__I0 (.I(\u_arbiter.i_wb_cpu_rdt[21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09081__I0 (.I(\u_arbiter.i_wb_cpu_rdt[22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08412__I0 (.I(\u_arbiter.i_wb_cpu_rdt[22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08223__A1 (.I(\u_arbiter.i_wb_cpu_rdt[22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05903__I0 (.I(\u_arbiter.i_wb_cpu_rdt[22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09083__I0 (.I(\u_arbiter.i_wb_cpu_rdt[23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08470__I0 (.I(\u_arbiter.i_wb_cpu_rdt[23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08226__A1 (.I(\u_arbiter.i_wb_cpu_rdt[23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05905__I0 (.I(\u_arbiter.i_wb_cpu_rdt[23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09085__I0 (.I(\u_arbiter.i_wb_cpu_rdt[24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08484__I0 (.I(\u_arbiter.i_wb_cpu_rdt[24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08229__A1 (.I(\u_arbiter.i_wb_cpu_rdt[24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05907__I0 (.I(\u_arbiter.i_wb_cpu_rdt[24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09087__I0 (.I(\u_arbiter.i_wb_cpu_rdt[25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08496__I0 (.I(\u_arbiter.i_wb_cpu_rdt[25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08232__A1 (.I(\u_arbiter.i_wb_cpu_rdt[25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05909__I0 (.I(\u_arbiter.i_wb_cpu_rdt[25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09089__I0 (.I(\u_arbiter.i_wb_cpu_rdt[26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08441__I0 (.I(\u_arbiter.i_wb_cpu_rdt[26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08234__A1 (.I(\u_arbiter.i_wb_cpu_rdt[26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05911__I0 (.I(\u_arbiter.i_wb_cpu_rdt[26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09091__A1 (.I(\u_arbiter.i_wb_cpu_rdt[27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08512__I0 (.I(\u_arbiter.i_wb_cpu_rdt[27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08237__A1 (.I(\u_arbiter.i_wb_cpu_rdt[27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05913__I0 (.I(\u_arbiter.i_wb_cpu_rdt[27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09093__I0 (.I(\u_arbiter.i_wb_cpu_rdt[28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08525__I0 (.I(\u_arbiter.i_wb_cpu_rdt[28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08240__A1 (.I(\u_arbiter.i_wb_cpu_rdt[28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05915__I0 (.I(\u_arbiter.i_wb_cpu_rdt[28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09095__I0 (.I(\u_arbiter.i_wb_cpu_rdt[29] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08532__I0 (.I(\u_arbiter.i_wb_cpu_rdt[29] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08242__A1 (.I(\u_arbiter.i_wb_cpu_rdt[29] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05918__A1 (.I(\u_arbiter.i_wb_cpu_rdt[29] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09097__I0 (.I(\u_arbiter.i_wb_cpu_rdt[30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08538__I0 (.I(\u_arbiter.i_wb_cpu_rdt[30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08244__A1 (.I(\u_arbiter.i_wb_cpu_rdt[30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05920__I0 (.I(\u_arbiter.i_wb_cpu_rdt[30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09099__I0 (.I(\u_arbiter.i_wb_cpu_rdt[31] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08643__I0 (.I(\u_arbiter.i_wb_cpu_rdt[31] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08246__A1 (.I(\u_arbiter.i_wb_cpu_rdt[31] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05922__I0 (.I(\u_arbiter.i_wb_cpu_rdt[31] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08390__I1 (.I(\u_arbiter.i_wb_cpu_rdt[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08332__A2 (.I(\u_arbiter.i_wb_cpu_rdt[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08317__I0 (.I(\u_arbiter.i_wb_cpu_rdt[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08167__A1 (.I(\u_arbiter.i_wb_cpu_rdt[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05866__I0 (.I(\u_arbiter.i_wb_cpu_rdt[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08401__I1 (.I(\u_arbiter.i_wb_cpu_rdt[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08355__A2 (.I(\u_arbiter.i_wb_cpu_rdt[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08313__I0 (.I(\u_arbiter.i_wb_cpu_rdt[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08169__A1 (.I(\u_arbiter.i_wb_cpu_rdt[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05868__I0 (.I(\u_arbiter.i_wb_cpu_rdt[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08412__I1 (.I(\u_arbiter.i_wb_cpu_rdt[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08312__I0 (.I(\u_arbiter.i_wb_cpu_rdt[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08175__A1 (.I(\u_arbiter.i_wb_cpu_rdt[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05870__I0 (.I(\u_arbiter.i_wb_cpu_rdt[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08470__I1 (.I(\u_arbiter.i_wb_cpu_rdt[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08297__I0 (.I(\u_arbiter.i_wb_cpu_rdt[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08178__A1 (.I(\u_arbiter.i_wb_cpu_rdt[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05872__I0 (.I(\u_arbiter.i_wb_cpu_rdt[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08484__I1 (.I(\u_arbiter.i_wb_cpu_rdt[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08304__I0 (.I(\u_arbiter.i_wb_cpu_rdt[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08300__A2 (.I(\u_arbiter.i_wb_cpu_rdt[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08181__A1 (.I(\u_arbiter.i_wb_cpu_rdt[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05874__I0 (.I(\u_arbiter.i_wb_cpu_rdt[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08496__I1 (.I(\u_arbiter.i_wb_cpu_rdt[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08296__I0 (.I(\u_arbiter.i_wb_cpu_rdt[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08184__A1 (.I(\u_arbiter.i_wb_cpu_rdt[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05876__I0 (.I(\u_arbiter.i_wb_cpu_rdt[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07856__A1 (.I(\u_cpu.cpu.alu.i_rs1 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06101__A1 (.I(\u_cpu.cpu.alu.i_rs1 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06096__A1 (.I(\u_cpu.cpu.alu.i_rs1 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05773__A1 (.I(\u_cpu.cpu.alu.i_rs1 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05771__A1 (.I(\u_cpu.cpu.alu.i_rs1 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05769__A1 (.I(\u_cpu.cpu.alu.i_rs1 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05708__A2 (.I(\u_cpu.cpu.alu.i_rs1 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05702__A1 (.I(\u_cpu.cpu.alu.i_rs1 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05685__A1 (.I(\u_cpu.cpu.alu.i_rs1 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07855__A1 (.I(\u_cpu.cpu.bne_or_bge ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05860__A1 (.I(\u_cpu.cpu.bne_or_bge ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05850__A1 (.I(\u_cpu.cpu.bne_or_bge ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05772__A1 (.I(\u_cpu.cpu.bne_or_bge ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05710__I (.I(\u_cpu.cpu.bne_or_bge ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05706__A2 (.I(\u_cpu.cpu.bne_or_bge ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05683__A2 (.I(\u_cpu.cpu.bne_or_bge ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04863__A2 (.I(\u_cpu.cpu.bne_or_bge ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04856__A2 (.I(\u_cpu.cpu.bne_or_bge ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09045__A1 (.I(\u_cpu.cpu.bufreg.i_sh_signed ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08750__A1 (.I(\u_cpu.cpu.bufreg.i_sh_signed ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05684__A2 (.I(\u_cpu.cpu.bufreg.i_sh_signed ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09524__A1 (.I(\u_cpu.cpu.ctrl.i_iscomp ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05787__A2 (.I(\u_cpu.cpu.ctrl.i_iscomp ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05786__A2 (.I(\u_cpu.cpu.ctrl.i_iscomp ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08812__A1 (.I(\u_cpu.cpu.ctrl.o_ibus_adr[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08810__B2 (.I(\u_cpu.cpu.ctrl.o_ibus_adr[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06015__A4 (.I(\u_cpu.cpu.ctrl.o_ibus_adr[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06009__A2 (.I(\u_cpu.cpu.ctrl.o_ibus_adr[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06005__A1 (.I(\u_cpu.cpu.ctrl.o_ibus_adr[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06002__A1 (.I(\u_cpu.cpu.ctrl.o_ibus_adr[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08798__A1 (.I(\u_cpu.cpu.ctrl.o_ibus_adr[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08796__B2 (.I(\u_cpu.cpu.ctrl.o_ibus_adr[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05973__A1 (.I(\u_cpu.cpu.ctrl.o_ibus_adr[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05969__A1 (.I(\u_cpu.cpu.ctrl.o_ibus_adr[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09515__A1 (.I(\u_cpu.cpu.decode.co_ebreak ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06125__A2 (.I(\u_cpu.cpu.decode.co_ebreak ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05750__I (.I(\u_cpu.cpu.decode.co_ebreak ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05721__A2 (.I(\u_cpu.cpu.decode.co_ebreak ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04889__A2 (.I(\u_cpu.cpu.decode.co_ebreak ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04862__B (.I(\u_cpu.cpu.decode.co_ebreak ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09492__A1 (.I(\u_cpu.cpu.decode.op21 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04872__A1 (.I(\u_cpu.cpu.decode.op21 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04868__A1 (.I(\u_cpu.cpu.decode.op21 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04861__I (.I(\u_cpu.cpu.decode.op21 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06125__A1 (.I(\u_cpu.cpu.decode.op26 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05717__A1 (.I(\u_cpu.cpu.decode.op26 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04889__A1 (.I(\u_cpu.cpu.decode.op26 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04867__I (.I(\u_cpu.cpu.decode.op26 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04862__A2 (.I(\u_cpu.cpu.decode.op26 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09099__I1 (.I(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08319__I1 (.I(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08279__A2 (.I(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09077__I1 (.I(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08331__A2 (.I(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08317__I1 (.I(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08649__A3 (.I(\u_cpu.cpu.genblk3.csr.i_mtip ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05845__A2 (.I(\u_cpu.cpu.genblk3.csr.i_mtip ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09522__A1 (.I(\u_cpu.cpu.genblk3.csr.mstatus_mie ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09512__A1 (.I(\u_cpu.cpu.genblk3.csr.mstatus_mie ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08649__A2 (.I(\u_cpu.cpu.genblk3.csr.mstatus_mie ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05724__B2 (.I(\u_cpu.cpu.genblk3.csr.mstatus_mie ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09526__A1 (.I(\u_cpu.cpu.genblk3.csr.o_new_irq ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09493__A1 (.I(\u_cpu.cpu.genblk3.csr.o_new_irq ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05732__A1 (.I(\u_cpu.cpu.genblk3.csr.o_new_irq ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04871__I (.I(\u_cpu.cpu.genblk3.csr.o_new_irq ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04864__B (.I(\u_cpu.cpu.genblk3.csr.o_new_irq ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08937__A1 (.I(\u_cpu.cpu.immdec.imm11_7[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08928__A1 (.I(\u_cpu.cpu.immdec.imm11_7[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06127__A1 (.I(\u_cpu.cpu.immdec.imm11_7[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06117__A1 (.I(\u_cpu.cpu.immdec.imm11_7[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08853__A1 (.I(\u_cpu.cpu.immdec.imm11_7[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06368__A1 (.I(\u_cpu.cpu.immdec.imm11_7[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06283__I (.I(\u_cpu.cpu.immdec.imm11_7[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06135__A1 (.I(\u_cpu.cpu.immdec.imm11_7[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06117__A2 (.I(\u_cpu.cpu.immdec.imm11_7[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08953__A1 (.I(\u_cpu.cpu.immdec.imm11_7[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08950__A1 (.I(\u_cpu.cpu.immdec.imm11_7[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06284__A1 (.I(\u_cpu.cpu.immdec.imm11_7[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06199__A1 (.I(\u_cpu.cpu.immdec.imm11_7[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06140__A1 (.I(\u_cpu.cpu.immdec.imm11_7[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06117__A3 (.I(\u_cpu.cpu.immdec.imm11_7[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08952__A1 (.I(\u_cpu.cpu.immdec.imm11_7[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06445__A2 (.I(\u_cpu.cpu.immdec.imm11_7[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06368__A2 (.I(\u_cpu.cpu.immdec.imm11_7[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06286__A1 (.I(\u_cpu.cpu.immdec.imm11_7[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06199__A2 (.I(\u_cpu.cpu.immdec.imm11_7[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06136__I (.I(\u_cpu.cpu.immdec.imm11_7[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06119__A1 (.I(\u_cpu.cpu.immdec.imm11_7[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08608__A1 (.I(\u_cpu.cpu.immdec.imm19_12_20[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08592__A1 (.I(\u_cpu.cpu.immdec.imm19_12_20[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04887__A1 (.I(\u_cpu.cpu.immdec.imm19_12_20[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08641__A1 (.I(\u_cpu.cpu.immdec.imm19_12_20[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08630__A1 (.I(\u_cpu.cpu.immdec.imm19_12_20[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04881__A1 (.I(\u_cpu.cpu.immdec.imm19_12_20[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08463__A1 (.I(\u_cpu.cpu.immdec.imm24_20[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05691__B (.I(\u_cpu.cpu.immdec.imm24_20[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04853__I (.I(\u_cpu.cpu.immdec.imm24_20[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08467__I (.I(\u_cpu.cpu.immdec.imm24_20[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08465__B2 (.I(\u_cpu.cpu.immdec.imm24_20[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04897__A1 (.I(\u_cpu.cpu.immdec.imm24_20[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08480__A1 (.I(\u_cpu.cpu.immdec.imm24_20[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08468__A1 (.I(\u_cpu.cpu.immdec.imm24_20[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04901__A1 (.I(\u_cpu.cpu.immdec.imm24_20[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08488__A1 (.I(\u_cpu.cpu.immdec.imm24_20[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08479__A1 (.I(\u_cpu.cpu.immdec.imm24_20[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04883__A1 (.I(\u_cpu.cpu.immdec.imm24_20[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08963__A1 (.I(\u_cpu.cpu.immdec.imm30_25[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08502__A1 (.I(\u_cpu.cpu.immdec.imm30_25[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08488__B2 (.I(\u_cpu.cpu.immdec.imm30_25[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08645__A1 (.I(\u_cpu.cpu.immdec.imm31 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05745__A1 (.I(\u_cpu.cpu.immdec.imm31 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05693__A2 (.I(\u_cpu.cpu.immdec.imm31 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09515__A2 (.I(\u_cpu.cpu.mem_bytecnt[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08132__A1 (.I(\u_cpu.cpu.mem_bytecnt[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08131__A1 (.I(\u_cpu.cpu.mem_bytecnt[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07867__A1 (.I(\u_cpu.cpu.mem_bytecnt[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07803__A1 (.I(\u_cpu.cpu.mem_bytecnt[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05779__A2 (.I(\u_cpu.cpu.mem_bytecnt[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05748__B (.I(\u_cpu.cpu.mem_bytecnt[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05716__A1 (.I(\u_cpu.cpu.mem_bytecnt[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11084__D (.I(\u_cpu.cpu.o_wdata1 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09498__B2 (.I(\u_cpu.cpu.state.genblk1.misalign_trap_sync_r ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09494__A1 (.I(\u_cpu.cpu.state.genblk1.misalign_trap_sync_r ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07852__A1 (.I(\u_cpu.cpu.state.genblk1.misalign_trap_sync_r ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06602__A1 (.I(\u_cpu.cpu.state.genblk1.misalign_trap_sync_r ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06587__A1 (.I(\u_cpu.cpu.state.genblk1.misalign_trap_sync_r ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05727__A1 (.I(\u_cpu.cpu.state.genblk1.misalign_trap_sync_r ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04873__A1 (.I(\u_cpu.cpu.state.genblk1.misalign_trap_sync_r ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04864__C (.I(\u_cpu.cpu.state.genblk1.misalign_trap_sync_r ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07869__A1 (.I(\u_cpu.cpu.state.init_done ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05833__A1 (.I(\u_cpu.cpu.state.init_done ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05740__C (.I(\u_cpu.cpu.state.init_done ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05732__A2 (.I(\u_cpu.cpu.state.init_done ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08754__A2 (.I(\u_cpu.cpu.state.o_cnt_r[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07810__A2 (.I(\u_cpu.cpu.state.o_cnt_r[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05832__A2 (.I(\u_cpu.cpu.state.o_cnt_r[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05759__A1 (.I(\u_cpu.cpu.state.o_cnt_r[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05681__A2 (.I(\u_cpu.cpu.state.o_cnt_r[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07808__A1 (.I(\u_cpu.cpu.state.o_cnt_r[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07798__A1 (.I(\u_cpu.cpu.state.o_cnt_r[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07797__A1 (.I(\u_cpu.cpu.state.o_cnt_r[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05832__A3 (.I(\u_cpu.cpu.state.o_cnt_r[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05718__A1 (.I(\u_cpu.cpu.state.o_cnt_r[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05681__A3 (.I(\u_cpu.cpu.state.o_cnt_r[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09606__A1 (.I(\u_cpu.rf_ram.memory[0][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05164__I0 (.I(\u_cpu.rf_ram.memory[0][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09608__A1 (.I(\u_cpu.rf_ram.memory[0][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05252__I0 (.I(\u_cpu.rf_ram.memory[0][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09612__A1 (.I(\u_cpu.rf_ram.memory[0][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05428__I0 (.I(\u_cpu.rf_ram.memory[0][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06676__A1 (.I(\u_cpu.rf_ram.memory[119][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05206__I3 (.I(\u_cpu.rf_ram.memory[119][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06678__A1 (.I(\u_cpu.rf_ram.memory[119][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05294__I3 (.I(\u_cpu.rf_ram.memory[119][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06680__A1 (.I(\u_cpu.rf_ram.memory[119][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05382__I3 (.I(\u_cpu.rf_ram.memory[119][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07634__A1 (.I(\u_cpu.rf_ram.memory[128][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05058__I0 (.I(\u_cpu.rf_ram.memory[128][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07636__A1 (.I(\u_cpu.rf_ram.memory[128][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05142__I0 (.I(\u_cpu.rf_ram.memory[128][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07640__A1 (.I(\u_cpu.rf_ram.memory[128][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05318__I0 (.I(\u_cpu.rf_ram.memory[128][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07642__A1 (.I(\u_cpu.rf_ram.memory[128][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05410__I0 (.I(\u_cpu.rf_ram.memory[128][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07646__A1 (.I(\u_cpu.rf_ram.memory[128][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05582__I0 (.I(\u_cpu.rf_ram.memory[128][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06709__A1 (.I(\u_cpu.rf_ram.memory[139][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05051__I3 (.I(\u_cpu.rf_ram.memory[139][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06711__A1 (.I(\u_cpu.rf_ram.memory[139][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05146__I3 (.I(\u_cpu.rf_ram.memory[139][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06713__A1 (.I(\u_cpu.rf_ram.memory[139][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05230__I3 (.I(\u_cpu.rf_ram.memory[139][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06715__A1 (.I(\u_cpu.rf_ram.memory[139][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05322__I3 (.I(\u_cpu.rf_ram.memory[139][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06721__A1 (.I(\u_cpu.rf_ram.memory[139][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05586__I3 (.I(\u_cpu.rf_ram.memory[139][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06723__A1 (.I(\u_cpu.rf_ram.memory[139][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05676__I3 (.I(\u_cpu.rf_ram.memory[139][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07010__A1 (.I(\u_cpu.rf_ram.memory[19][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05159__I3 (.I(\u_cpu.rf_ram.memory[19][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07020__A1 (.I(\u_cpu.rf_ram.memory[19][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05599__I3 (.I(\u_cpu.rf_ram.memory[19][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07609__A1 (.I(\u_cpu.rf_ram.memory[22][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04929__I2 (.I(\u_cpu.rf_ram.memory[22][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07612__A1 (.I(\u_cpu.rf_ram.memory[22][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05069__I2 (.I(\u_cpu.rf_ram.memory[22][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07618__A1 (.I(\u_cpu.rf_ram.memory[22][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05245__I2 (.I(\u_cpu.rf_ram.memory[22][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07621__A1 (.I(\u_cpu.rf_ram.memory[22][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05333__I2 (.I(\u_cpu.rf_ram.memory[22][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07624__A1 (.I(\u_cpu.rf_ram.memory[22][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05421__I2 (.I(\u_cpu.rf_ram.memory[22][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07627__A1 (.I(\u_cpu.rf_ram.memory[22][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05509__I2 (.I(\u_cpu.rf_ram.memory[22][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07630__A1 (.I(\u_cpu.rf_ram.memory[22][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05597__I2 (.I(\u_cpu.rf_ram.memory[22][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08904__A1 (.I(\u_cpu.rf_ram.memory[2][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05516__I2 (.I(\u_cpu.rf_ram.memory[2][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07446__A1 (.I(\u_cpu.rf_ram.memory[49][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04993__I1 (.I(\u_cpu.rf_ram.memory[49][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07448__A1 (.I(\u_cpu.rf_ram.memory[49][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05098__I1 (.I(\u_cpu.rf_ram.memory[49][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07452__A1 (.I(\u_cpu.rf_ram.memory[49][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05274__I1 (.I(\u_cpu.rf_ram.memory[49][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07454__A1 (.I(\u_cpu.rf_ram.memory[49][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05362__I1 (.I(\u_cpu.rf_ram.memory[49][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07456__A1 (.I(\u_cpu.rf_ram.memory[49][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05450__I1 (.I(\u_cpu.rf_ram.memory[49][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07458__A1 (.I(\u_cpu.rf_ram.memory[49][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05538__I1 (.I(\u_cpu.rf_ram.memory[49][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06172__A1 (.I(\u_cpu.rf_ram.memory[82][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05390__I2 (.I(\u_cpu.rf_ram.memory[82][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06178__A1 (.I(\u_cpu.rf_ram.memory[82][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05478__I2 (.I(\u_cpu.rf_ram.memory[82][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06184__A1 (.I(\u_cpu.rf_ram.memory[82][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05566__I2 (.I(\u_cpu.rf_ram.memory[82][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06190__A1 (.I(\u_cpu.rf_ram.memory[82][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05654__I2 (.I(\u_cpu.rf_ram.memory[82][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11075__D (.I(\u_cpu.rf_ram_if.rtrig0 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09695__A3 (.I(\u_cpu.rf_ram_if.rtrig0 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06137__B1 (.I(\u_cpu.rf_ram_if.rtrig0 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04919__A2 (.I(\u_cpu.rf_ram_if.rtrig0 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04887__A2 (.I(\u_cpu.rf_ram_if.rtrig0 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04879__A1 (.I(\u_cpu.rf_ram_if.rtrig0 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04874__B (.I(\u_cpu.rf_ram_if.rtrig0 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11069__D (.I(\u_cpu.rf_ram_if.wdata0_r[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06181__A2 (.I(\u_cpu.rf_ram_if.wdata0_r[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11083__D (.I(\u_cpu.rf_ram_if.wdata1_r[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06186__I (.I(\u_cpu.rf_ram_if.wdata1_r[7] ));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_1_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_1_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_3_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_3_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_4_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_4_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_4_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_6_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_6_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_9_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_10_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_10_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_10_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_13_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_14_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_15_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_16_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_17_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_18_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_20_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_21_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_22_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_22_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_23_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_24_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_24_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_25_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_26_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_26_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_28_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_32_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_34_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_36_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_36_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_35 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_37_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_38_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_35 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_39_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_40_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_40_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_41_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_41_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_41_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_11 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_44_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_44_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_45_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_46_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_47_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_48_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_48_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_48_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_49_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_50_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_51_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_52_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_53_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_54_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_55_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_55_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_56_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_57_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_11 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_58_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_59_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_59_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_60_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_62_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_62_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_63_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_64_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_66_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_68_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_69_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_70_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_71_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_72_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_76_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_77_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_80_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_80_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_11 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_82_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_84_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_35 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_88_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_88_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_96_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_98_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_100_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_104_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_106_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_108_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_110_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_113_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_114_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_114_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_114_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_115_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_116_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_116_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_116_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_118_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_118_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_119_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_120_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_120_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_120_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_121_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_122_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_122_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_124_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_124_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_124_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_126_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_126_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_126_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_127_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_128_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_128_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_129_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_129_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_131_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_131_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_132_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_132_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_133_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_133_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_134_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_134_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_134_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_136_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_136_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_137_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_137_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_138_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_138_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_138_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_138_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_138_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_139_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_139_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_139_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_139_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_140_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_140_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_140_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_140_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_140_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_141_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_141_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_141_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_141_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_141_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_142_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_142_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_142_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_142_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_142_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_142_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_142_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_142_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_142_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_143_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_143_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_143_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_143_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_1192 ();
endmodule

