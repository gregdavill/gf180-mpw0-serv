// This is the unpowered netlist.
module serv_1 (io_in,
    io_oeb,
    io_out);
 input [4:0] io_in;
 output [4:0] io_oeb;
 output [4:0] io_out;

 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire _04725_;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire _04785_;
 wire _04786_;
 wire _04787_;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire _04809_;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire _04818_;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire \u_arbiter.i_wb_cpu_ack ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[10] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[11] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[12] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[13] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[14] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[15] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[16] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[17] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[18] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[19] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[20] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[21] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[22] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[23] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[24] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[25] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[26] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[27] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[28] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[29] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[2] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[30] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[31] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[3] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[4] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[5] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[6] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[7] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[8] ;
 wire \u_arbiter.i_wb_cpu_dbus_adr[9] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[0] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[10] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[11] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[12] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[13] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[14] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[15] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[16] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[17] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[18] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[19] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[1] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[20] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[21] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[22] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[23] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[24] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[25] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[26] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[27] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[28] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[29] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[2] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[30] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[31] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[3] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[4] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[5] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[6] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[7] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[8] ;
 wire \u_arbiter.i_wb_cpu_dbus_dat[9] ;
 wire \u_arbiter.i_wb_cpu_dbus_sel[0] ;
 wire \u_arbiter.i_wb_cpu_dbus_sel[1] ;
 wire \u_arbiter.i_wb_cpu_dbus_sel[2] ;
 wire \u_arbiter.i_wb_cpu_dbus_sel[3] ;
 wire \u_arbiter.i_wb_cpu_dbus_we ;
 wire \u_arbiter.i_wb_cpu_ibus_adr[0] ;
 wire \u_arbiter.i_wb_cpu_ibus_adr[1] ;
 wire \u_arbiter.i_wb_cpu_rdt[0] ;
 wire \u_arbiter.i_wb_cpu_rdt[10] ;
 wire \u_arbiter.i_wb_cpu_rdt[11] ;
 wire \u_arbiter.i_wb_cpu_rdt[12] ;
 wire \u_arbiter.i_wb_cpu_rdt[13] ;
 wire \u_arbiter.i_wb_cpu_rdt[14] ;
 wire \u_arbiter.i_wb_cpu_rdt[15] ;
 wire \u_arbiter.i_wb_cpu_rdt[16] ;
 wire \u_arbiter.i_wb_cpu_rdt[17] ;
 wire \u_arbiter.i_wb_cpu_rdt[18] ;
 wire \u_arbiter.i_wb_cpu_rdt[19] ;
 wire \u_arbiter.i_wb_cpu_rdt[1] ;
 wire \u_arbiter.i_wb_cpu_rdt[20] ;
 wire \u_arbiter.i_wb_cpu_rdt[21] ;
 wire \u_arbiter.i_wb_cpu_rdt[22] ;
 wire \u_arbiter.i_wb_cpu_rdt[23] ;
 wire \u_arbiter.i_wb_cpu_rdt[24] ;
 wire \u_arbiter.i_wb_cpu_rdt[25] ;
 wire \u_arbiter.i_wb_cpu_rdt[26] ;
 wire \u_arbiter.i_wb_cpu_rdt[27] ;
 wire \u_arbiter.i_wb_cpu_rdt[28] ;
 wire \u_arbiter.i_wb_cpu_rdt[29] ;
 wire \u_arbiter.i_wb_cpu_rdt[2] ;
 wire \u_arbiter.i_wb_cpu_rdt[30] ;
 wire \u_arbiter.i_wb_cpu_rdt[31] ;
 wire \u_arbiter.i_wb_cpu_rdt[3] ;
 wire \u_arbiter.i_wb_cpu_rdt[4] ;
 wire \u_arbiter.i_wb_cpu_rdt[5] ;
 wire \u_arbiter.i_wb_cpu_rdt[6] ;
 wire \u_arbiter.i_wb_cpu_rdt[7] ;
 wire \u_arbiter.i_wb_cpu_rdt[8] ;
 wire \u_arbiter.i_wb_cpu_rdt[9] ;
 wire \u_arbiter.o_wb_cpu_adr[0] ;
 wire \u_arbiter.o_wb_cpu_adr[10] ;
 wire \u_arbiter.o_wb_cpu_adr[11] ;
 wire \u_arbiter.o_wb_cpu_adr[12] ;
 wire \u_arbiter.o_wb_cpu_adr[13] ;
 wire \u_arbiter.o_wb_cpu_adr[14] ;
 wire \u_arbiter.o_wb_cpu_adr[15] ;
 wire \u_arbiter.o_wb_cpu_adr[16] ;
 wire \u_arbiter.o_wb_cpu_adr[17] ;
 wire \u_arbiter.o_wb_cpu_adr[18] ;
 wire \u_arbiter.o_wb_cpu_adr[19] ;
 wire \u_arbiter.o_wb_cpu_adr[1] ;
 wire \u_arbiter.o_wb_cpu_adr[20] ;
 wire \u_arbiter.o_wb_cpu_adr[21] ;
 wire \u_arbiter.o_wb_cpu_adr[22] ;
 wire \u_arbiter.o_wb_cpu_adr[23] ;
 wire \u_arbiter.o_wb_cpu_adr[24] ;
 wire \u_arbiter.o_wb_cpu_adr[25] ;
 wire \u_arbiter.o_wb_cpu_adr[26] ;
 wire \u_arbiter.o_wb_cpu_adr[27] ;
 wire \u_arbiter.o_wb_cpu_adr[28] ;
 wire \u_arbiter.o_wb_cpu_adr[29] ;
 wire \u_arbiter.o_wb_cpu_adr[2] ;
 wire \u_arbiter.o_wb_cpu_adr[30] ;
 wire \u_arbiter.o_wb_cpu_adr[31] ;
 wire \u_arbiter.o_wb_cpu_adr[3] ;
 wire \u_arbiter.o_wb_cpu_adr[4] ;
 wire \u_arbiter.o_wb_cpu_adr[5] ;
 wire \u_arbiter.o_wb_cpu_adr[6] ;
 wire \u_arbiter.o_wb_cpu_adr[7] ;
 wire \u_arbiter.o_wb_cpu_adr[8] ;
 wire \u_arbiter.o_wb_cpu_adr[9] ;
 wire \u_arbiter.o_wb_cpu_cyc ;
 wire \u_arbiter.o_wb_cpu_we ;
 wire \u_cpu.cpu.alu.add_cy_r ;
 wire \u_cpu.cpu.alu.cmp_r ;
 wire \u_cpu.cpu.alu.i_rs1 ;
 wire \u_cpu.cpu.bne_or_bge ;
 wire \u_cpu.cpu.branch_op ;
 wire \u_cpu.cpu.bufreg.c_r ;
 wire \u_cpu.cpu.bufreg.i_sh_signed ;
 wire \u_cpu.cpu.bufreg.lsb[0] ;
 wire \u_cpu.cpu.bufreg.lsb[1] ;
 wire \u_cpu.cpu.bufreg2.i_cnt_done ;
 wire \u_cpu.cpu.csr_d_sel ;
 wire \u_cpu.cpu.csr_imm ;
 wire \u_cpu.cpu.ctrl.i_iscomp ;
 wire \u_cpu.cpu.ctrl.i_jump ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[10] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[11] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[12] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[13] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[14] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[15] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[16] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[17] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[18] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[19] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[20] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[21] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[22] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[23] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[24] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[25] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[26] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[27] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[28] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[29] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[2] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[30] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[31] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[3] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[4] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[5] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[6] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[7] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[8] ;
 wire \u_cpu.cpu.ctrl.o_ibus_adr[9] ;
 wire \u_cpu.cpu.ctrl.pc_plus_4_cy_r ;
 wire \u_cpu.cpu.ctrl.pc_plus_offset_cy_r ;
 wire \u_cpu.cpu.decode.co_ebreak ;
 wire \u_cpu.cpu.decode.co_mem_word ;
 wire \u_cpu.cpu.decode.op21 ;
 wire \u_cpu.cpu.decode.op22 ;
 wire \u_cpu.cpu.decode.op26 ;
 wire \u_cpu.cpu.decode.opcode[0] ;
 wire \u_cpu.cpu.decode.opcode[1] ;
 wire \u_cpu.cpu.decode.opcode[2] ;
 wire \u_cpu.cpu.genblk1.align.ctrl_misal ;
 wire \u_cpu.cpu.genblk1.align.ibus_rdt_concat[0] ;
 wire \u_cpu.cpu.genblk1.align.ibus_rdt_concat[10] ;
 wire \u_cpu.cpu.genblk1.align.ibus_rdt_concat[11] ;
 wire \u_cpu.cpu.genblk1.align.ibus_rdt_concat[12] ;
 wire \u_cpu.cpu.genblk1.align.ibus_rdt_concat[13] ;
 wire \u_cpu.cpu.genblk1.align.ibus_rdt_concat[14] ;
 wire \u_cpu.cpu.genblk1.align.ibus_rdt_concat[15] ;
 wire \u_cpu.cpu.genblk1.align.ibus_rdt_concat[1] ;
 wire \u_cpu.cpu.genblk1.align.ibus_rdt_concat[2] ;
 wire \u_cpu.cpu.genblk1.align.ibus_rdt_concat[3] ;
 wire \u_cpu.cpu.genblk1.align.ibus_rdt_concat[4] ;
 wire \u_cpu.cpu.genblk1.align.ibus_rdt_concat[5] ;
 wire \u_cpu.cpu.genblk1.align.ibus_rdt_concat[6] ;
 wire \u_cpu.cpu.genblk1.align.ibus_rdt_concat[7] ;
 wire \u_cpu.cpu.genblk1.align.ibus_rdt_concat[8] ;
 wire \u_cpu.cpu.genblk1.align.ibus_rdt_concat[9] ;
 wire \u_cpu.cpu.genblk3.csr.i_mtip ;
 wire \u_cpu.cpu.genblk3.csr.mcause31 ;
 wire \u_cpu.cpu.genblk3.csr.mcause3_0[0] ;
 wire \u_cpu.cpu.genblk3.csr.mcause3_0[1] ;
 wire \u_cpu.cpu.genblk3.csr.mcause3_0[2] ;
 wire \u_cpu.cpu.genblk3.csr.mcause3_0[3] ;
 wire \u_cpu.cpu.genblk3.csr.mie_mtie ;
 wire \u_cpu.cpu.genblk3.csr.mstatus_mie ;
 wire \u_cpu.cpu.genblk3.csr.mstatus_mpie ;
 wire \u_cpu.cpu.genblk3.csr.o_new_irq ;
 wire \u_cpu.cpu.genblk3.csr.timer_irq_r ;
 wire \u_cpu.cpu.immdec.imm11_7[0] ;
 wire \u_cpu.cpu.immdec.imm11_7[1] ;
 wire \u_cpu.cpu.immdec.imm11_7[2] ;
 wire \u_cpu.cpu.immdec.imm11_7[3] ;
 wire \u_cpu.cpu.immdec.imm11_7[4] ;
 wire \u_cpu.cpu.immdec.imm19_12_20[0] ;
 wire \u_cpu.cpu.immdec.imm19_12_20[1] ;
 wire \u_cpu.cpu.immdec.imm19_12_20[2] ;
 wire \u_cpu.cpu.immdec.imm19_12_20[3] ;
 wire \u_cpu.cpu.immdec.imm19_12_20[5] ;
 wire \u_cpu.cpu.immdec.imm19_12_20[6] ;
 wire \u_cpu.cpu.immdec.imm19_12_20[7] ;
 wire \u_cpu.cpu.immdec.imm19_12_20[8] ;
 wire \u_cpu.cpu.immdec.imm24_20[0] ;
 wire \u_cpu.cpu.immdec.imm24_20[1] ;
 wire \u_cpu.cpu.immdec.imm24_20[2] ;
 wire \u_cpu.cpu.immdec.imm24_20[3] ;
 wire \u_cpu.cpu.immdec.imm24_20[4] ;
 wire \u_cpu.cpu.immdec.imm30_25[0] ;
 wire \u_cpu.cpu.immdec.imm30_25[1] ;
 wire \u_cpu.cpu.immdec.imm30_25[2] ;
 wire \u_cpu.cpu.immdec.imm30_25[3] ;
 wire \u_cpu.cpu.immdec.imm30_25[4] ;
 wire \u_cpu.cpu.immdec.imm30_25[5] ;
 wire \u_cpu.cpu.immdec.imm31 ;
 wire \u_cpu.cpu.immdec.imm7 ;
 wire \u_cpu.cpu.mem_bytecnt[0] ;
 wire \u_cpu.cpu.mem_bytecnt[1] ;
 wire \u_cpu.cpu.mem_if.signbit ;
 wire \u_cpu.cpu.o_wdata0 ;
 wire \u_cpu.cpu.o_wdata1 ;
 wire \u_cpu.cpu.o_wen0 ;
 wire \u_cpu.cpu.o_wen1 ;
 wire \u_cpu.cpu.state.genblk1.misalign_trap_sync_r ;
 wire \u_cpu.cpu.state.ibus_cyc ;
 wire \u_cpu.cpu.state.init_done ;
 wire \u_cpu.cpu.state.o_cnt[2] ;
 wire \u_cpu.cpu.state.o_cnt_r[0] ;
 wire \u_cpu.cpu.state.o_cnt_r[1] ;
 wire \u_cpu.cpu.state.o_cnt_r[2] ;
 wire \u_cpu.cpu.state.o_cnt_r[3] ;
 wire \u_cpu.cpu.state.stage_two_req ;
 wire \u_cpu.raddr[0] ;
 wire \u_cpu.raddr[1] ;
 wire \u_cpu.rf_ram.memory[0][0] ;
 wire \u_cpu.rf_ram.memory[0][1] ;
 wire \u_cpu.rf_ram.memory[0][2] ;
 wire \u_cpu.rf_ram.memory[0][3] ;
 wire \u_cpu.rf_ram.memory[0][4] ;
 wire \u_cpu.rf_ram.memory[0][5] ;
 wire \u_cpu.rf_ram.memory[0][6] ;
 wire \u_cpu.rf_ram.memory[0][7] ;
 wire \u_cpu.rf_ram.memory[100][0] ;
 wire \u_cpu.rf_ram.memory[100][1] ;
 wire \u_cpu.rf_ram.memory[100][2] ;
 wire \u_cpu.rf_ram.memory[100][3] ;
 wire \u_cpu.rf_ram.memory[100][4] ;
 wire \u_cpu.rf_ram.memory[100][5] ;
 wire \u_cpu.rf_ram.memory[100][6] ;
 wire \u_cpu.rf_ram.memory[100][7] ;
 wire \u_cpu.rf_ram.memory[101][0] ;
 wire \u_cpu.rf_ram.memory[101][1] ;
 wire \u_cpu.rf_ram.memory[101][2] ;
 wire \u_cpu.rf_ram.memory[101][3] ;
 wire \u_cpu.rf_ram.memory[101][4] ;
 wire \u_cpu.rf_ram.memory[101][5] ;
 wire \u_cpu.rf_ram.memory[101][6] ;
 wire \u_cpu.rf_ram.memory[101][7] ;
 wire \u_cpu.rf_ram.memory[102][0] ;
 wire \u_cpu.rf_ram.memory[102][1] ;
 wire \u_cpu.rf_ram.memory[102][2] ;
 wire \u_cpu.rf_ram.memory[102][3] ;
 wire \u_cpu.rf_ram.memory[102][4] ;
 wire \u_cpu.rf_ram.memory[102][5] ;
 wire \u_cpu.rf_ram.memory[102][6] ;
 wire \u_cpu.rf_ram.memory[102][7] ;
 wire \u_cpu.rf_ram.memory[103][0] ;
 wire \u_cpu.rf_ram.memory[103][1] ;
 wire \u_cpu.rf_ram.memory[103][2] ;
 wire \u_cpu.rf_ram.memory[103][3] ;
 wire \u_cpu.rf_ram.memory[103][4] ;
 wire \u_cpu.rf_ram.memory[103][5] ;
 wire \u_cpu.rf_ram.memory[103][6] ;
 wire \u_cpu.rf_ram.memory[103][7] ;
 wire \u_cpu.rf_ram.memory[104][0] ;
 wire \u_cpu.rf_ram.memory[104][1] ;
 wire \u_cpu.rf_ram.memory[104][2] ;
 wire \u_cpu.rf_ram.memory[104][3] ;
 wire \u_cpu.rf_ram.memory[104][4] ;
 wire \u_cpu.rf_ram.memory[104][5] ;
 wire \u_cpu.rf_ram.memory[104][6] ;
 wire \u_cpu.rf_ram.memory[104][7] ;
 wire \u_cpu.rf_ram.memory[105][0] ;
 wire \u_cpu.rf_ram.memory[105][1] ;
 wire \u_cpu.rf_ram.memory[105][2] ;
 wire \u_cpu.rf_ram.memory[105][3] ;
 wire \u_cpu.rf_ram.memory[105][4] ;
 wire \u_cpu.rf_ram.memory[105][5] ;
 wire \u_cpu.rf_ram.memory[105][6] ;
 wire \u_cpu.rf_ram.memory[105][7] ;
 wire \u_cpu.rf_ram.memory[106][0] ;
 wire \u_cpu.rf_ram.memory[106][1] ;
 wire \u_cpu.rf_ram.memory[106][2] ;
 wire \u_cpu.rf_ram.memory[106][3] ;
 wire \u_cpu.rf_ram.memory[106][4] ;
 wire \u_cpu.rf_ram.memory[106][5] ;
 wire \u_cpu.rf_ram.memory[106][6] ;
 wire \u_cpu.rf_ram.memory[106][7] ;
 wire \u_cpu.rf_ram.memory[107][0] ;
 wire \u_cpu.rf_ram.memory[107][1] ;
 wire \u_cpu.rf_ram.memory[107][2] ;
 wire \u_cpu.rf_ram.memory[107][3] ;
 wire \u_cpu.rf_ram.memory[107][4] ;
 wire \u_cpu.rf_ram.memory[107][5] ;
 wire \u_cpu.rf_ram.memory[107][6] ;
 wire \u_cpu.rf_ram.memory[107][7] ;
 wire \u_cpu.rf_ram.memory[108][0] ;
 wire \u_cpu.rf_ram.memory[108][1] ;
 wire \u_cpu.rf_ram.memory[108][2] ;
 wire \u_cpu.rf_ram.memory[108][3] ;
 wire \u_cpu.rf_ram.memory[108][4] ;
 wire \u_cpu.rf_ram.memory[108][5] ;
 wire \u_cpu.rf_ram.memory[108][6] ;
 wire \u_cpu.rf_ram.memory[108][7] ;
 wire \u_cpu.rf_ram.memory[109][0] ;
 wire \u_cpu.rf_ram.memory[109][1] ;
 wire \u_cpu.rf_ram.memory[109][2] ;
 wire \u_cpu.rf_ram.memory[109][3] ;
 wire \u_cpu.rf_ram.memory[109][4] ;
 wire \u_cpu.rf_ram.memory[109][5] ;
 wire \u_cpu.rf_ram.memory[109][6] ;
 wire \u_cpu.rf_ram.memory[109][7] ;
 wire \u_cpu.rf_ram.memory[10][0] ;
 wire \u_cpu.rf_ram.memory[10][1] ;
 wire \u_cpu.rf_ram.memory[10][2] ;
 wire \u_cpu.rf_ram.memory[10][3] ;
 wire \u_cpu.rf_ram.memory[10][4] ;
 wire \u_cpu.rf_ram.memory[10][5] ;
 wire \u_cpu.rf_ram.memory[10][6] ;
 wire \u_cpu.rf_ram.memory[10][7] ;
 wire \u_cpu.rf_ram.memory[110][0] ;
 wire \u_cpu.rf_ram.memory[110][1] ;
 wire \u_cpu.rf_ram.memory[110][2] ;
 wire \u_cpu.rf_ram.memory[110][3] ;
 wire \u_cpu.rf_ram.memory[110][4] ;
 wire \u_cpu.rf_ram.memory[110][5] ;
 wire \u_cpu.rf_ram.memory[110][6] ;
 wire \u_cpu.rf_ram.memory[110][7] ;
 wire \u_cpu.rf_ram.memory[111][0] ;
 wire \u_cpu.rf_ram.memory[111][1] ;
 wire \u_cpu.rf_ram.memory[111][2] ;
 wire \u_cpu.rf_ram.memory[111][3] ;
 wire \u_cpu.rf_ram.memory[111][4] ;
 wire \u_cpu.rf_ram.memory[111][5] ;
 wire \u_cpu.rf_ram.memory[111][6] ;
 wire \u_cpu.rf_ram.memory[111][7] ;
 wire \u_cpu.rf_ram.memory[112][0] ;
 wire \u_cpu.rf_ram.memory[112][1] ;
 wire \u_cpu.rf_ram.memory[112][2] ;
 wire \u_cpu.rf_ram.memory[112][3] ;
 wire \u_cpu.rf_ram.memory[112][4] ;
 wire \u_cpu.rf_ram.memory[112][5] ;
 wire \u_cpu.rf_ram.memory[112][6] ;
 wire \u_cpu.rf_ram.memory[112][7] ;
 wire \u_cpu.rf_ram.memory[113][0] ;
 wire \u_cpu.rf_ram.memory[113][1] ;
 wire \u_cpu.rf_ram.memory[113][2] ;
 wire \u_cpu.rf_ram.memory[113][3] ;
 wire \u_cpu.rf_ram.memory[113][4] ;
 wire \u_cpu.rf_ram.memory[113][5] ;
 wire \u_cpu.rf_ram.memory[113][6] ;
 wire \u_cpu.rf_ram.memory[113][7] ;
 wire \u_cpu.rf_ram.memory[114][0] ;
 wire \u_cpu.rf_ram.memory[114][1] ;
 wire \u_cpu.rf_ram.memory[114][2] ;
 wire \u_cpu.rf_ram.memory[114][3] ;
 wire \u_cpu.rf_ram.memory[114][4] ;
 wire \u_cpu.rf_ram.memory[114][5] ;
 wire \u_cpu.rf_ram.memory[114][6] ;
 wire \u_cpu.rf_ram.memory[114][7] ;
 wire \u_cpu.rf_ram.memory[115][0] ;
 wire \u_cpu.rf_ram.memory[115][1] ;
 wire \u_cpu.rf_ram.memory[115][2] ;
 wire \u_cpu.rf_ram.memory[115][3] ;
 wire \u_cpu.rf_ram.memory[115][4] ;
 wire \u_cpu.rf_ram.memory[115][5] ;
 wire \u_cpu.rf_ram.memory[115][6] ;
 wire \u_cpu.rf_ram.memory[115][7] ;
 wire \u_cpu.rf_ram.memory[116][0] ;
 wire \u_cpu.rf_ram.memory[116][1] ;
 wire \u_cpu.rf_ram.memory[116][2] ;
 wire \u_cpu.rf_ram.memory[116][3] ;
 wire \u_cpu.rf_ram.memory[116][4] ;
 wire \u_cpu.rf_ram.memory[116][5] ;
 wire \u_cpu.rf_ram.memory[116][6] ;
 wire \u_cpu.rf_ram.memory[116][7] ;
 wire \u_cpu.rf_ram.memory[117][0] ;
 wire \u_cpu.rf_ram.memory[117][1] ;
 wire \u_cpu.rf_ram.memory[117][2] ;
 wire \u_cpu.rf_ram.memory[117][3] ;
 wire \u_cpu.rf_ram.memory[117][4] ;
 wire \u_cpu.rf_ram.memory[117][5] ;
 wire \u_cpu.rf_ram.memory[117][6] ;
 wire \u_cpu.rf_ram.memory[117][7] ;
 wire \u_cpu.rf_ram.memory[118][0] ;
 wire \u_cpu.rf_ram.memory[118][1] ;
 wire \u_cpu.rf_ram.memory[118][2] ;
 wire \u_cpu.rf_ram.memory[118][3] ;
 wire \u_cpu.rf_ram.memory[118][4] ;
 wire \u_cpu.rf_ram.memory[118][5] ;
 wire \u_cpu.rf_ram.memory[118][6] ;
 wire \u_cpu.rf_ram.memory[118][7] ;
 wire \u_cpu.rf_ram.memory[119][0] ;
 wire \u_cpu.rf_ram.memory[119][1] ;
 wire \u_cpu.rf_ram.memory[119][2] ;
 wire \u_cpu.rf_ram.memory[119][3] ;
 wire \u_cpu.rf_ram.memory[119][4] ;
 wire \u_cpu.rf_ram.memory[119][5] ;
 wire \u_cpu.rf_ram.memory[119][6] ;
 wire \u_cpu.rf_ram.memory[119][7] ;
 wire \u_cpu.rf_ram.memory[11][0] ;
 wire \u_cpu.rf_ram.memory[11][1] ;
 wire \u_cpu.rf_ram.memory[11][2] ;
 wire \u_cpu.rf_ram.memory[11][3] ;
 wire \u_cpu.rf_ram.memory[11][4] ;
 wire \u_cpu.rf_ram.memory[11][5] ;
 wire \u_cpu.rf_ram.memory[11][6] ;
 wire \u_cpu.rf_ram.memory[11][7] ;
 wire \u_cpu.rf_ram.memory[120][0] ;
 wire \u_cpu.rf_ram.memory[120][1] ;
 wire \u_cpu.rf_ram.memory[120][2] ;
 wire \u_cpu.rf_ram.memory[120][3] ;
 wire \u_cpu.rf_ram.memory[120][4] ;
 wire \u_cpu.rf_ram.memory[120][5] ;
 wire \u_cpu.rf_ram.memory[120][6] ;
 wire \u_cpu.rf_ram.memory[120][7] ;
 wire \u_cpu.rf_ram.memory[121][0] ;
 wire \u_cpu.rf_ram.memory[121][1] ;
 wire \u_cpu.rf_ram.memory[121][2] ;
 wire \u_cpu.rf_ram.memory[121][3] ;
 wire \u_cpu.rf_ram.memory[121][4] ;
 wire \u_cpu.rf_ram.memory[121][5] ;
 wire \u_cpu.rf_ram.memory[121][6] ;
 wire \u_cpu.rf_ram.memory[121][7] ;
 wire \u_cpu.rf_ram.memory[122][0] ;
 wire \u_cpu.rf_ram.memory[122][1] ;
 wire \u_cpu.rf_ram.memory[122][2] ;
 wire \u_cpu.rf_ram.memory[122][3] ;
 wire \u_cpu.rf_ram.memory[122][4] ;
 wire \u_cpu.rf_ram.memory[122][5] ;
 wire \u_cpu.rf_ram.memory[122][6] ;
 wire \u_cpu.rf_ram.memory[122][7] ;
 wire \u_cpu.rf_ram.memory[123][0] ;
 wire \u_cpu.rf_ram.memory[123][1] ;
 wire \u_cpu.rf_ram.memory[123][2] ;
 wire \u_cpu.rf_ram.memory[123][3] ;
 wire \u_cpu.rf_ram.memory[123][4] ;
 wire \u_cpu.rf_ram.memory[123][5] ;
 wire \u_cpu.rf_ram.memory[123][6] ;
 wire \u_cpu.rf_ram.memory[123][7] ;
 wire \u_cpu.rf_ram.memory[124][0] ;
 wire \u_cpu.rf_ram.memory[124][1] ;
 wire \u_cpu.rf_ram.memory[124][2] ;
 wire \u_cpu.rf_ram.memory[124][3] ;
 wire \u_cpu.rf_ram.memory[124][4] ;
 wire \u_cpu.rf_ram.memory[124][5] ;
 wire \u_cpu.rf_ram.memory[124][6] ;
 wire \u_cpu.rf_ram.memory[124][7] ;
 wire \u_cpu.rf_ram.memory[125][0] ;
 wire \u_cpu.rf_ram.memory[125][1] ;
 wire \u_cpu.rf_ram.memory[125][2] ;
 wire \u_cpu.rf_ram.memory[125][3] ;
 wire \u_cpu.rf_ram.memory[125][4] ;
 wire \u_cpu.rf_ram.memory[125][5] ;
 wire \u_cpu.rf_ram.memory[125][6] ;
 wire \u_cpu.rf_ram.memory[125][7] ;
 wire \u_cpu.rf_ram.memory[126][0] ;
 wire \u_cpu.rf_ram.memory[126][1] ;
 wire \u_cpu.rf_ram.memory[126][2] ;
 wire \u_cpu.rf_ram.memory[126][3] ;
 wire \u_cpu.rf_ram.memory[126][4] ;
 wire \u_cpu.rf_ram.memory[126][5] ;
 wire \u_cpu.rf_ram.memory[126][6] ;
 wire \u_cpu.rf_ram.memory[126][7] ;
 wire \u_cpu.rf_ram.memory[127][0] ;
 wire \u_cpu.rf_ram.memory[127][1] ;
 wire \u_cpu.rf_ram.memory[127][2] ;
 wire \u_cpu.rf_ram.memory[127][3] ;
 wire \u_cpu.rf_ram.memory[127][4] ;
 wire \u_cpu.rf_ram.memory[127][5] ;
 wire \u_cpu.rf_ram.memory[127][6] ;
 wire \u_cpu.rf_ram.memory[127][7] ;
 wire \u_cpu.rf_ram.memory[128][0] ;
 wire \u_cpu.rf_ram.memory[128][1] ;
 wire \u_cpu.rf_ram.memory[128][2] ;
 wire \u_cpu.rf_ram.memory[128][3] ;
 wire \u_cpu.rf_ram.memory[128][4] ;
 wire \u_cpu.rf_ram.memory[128][5] ;
 wire \u_cpu.rf_ram.memory[128][6] ;
 wire \u_cpu.rf_ram.memory[128][7] ;
 wire \u_cpu.rf_ram.memory[129][0] ;
 wire \u_cpu.rf_ram.memory[129][1] ;
 wire \u_cpu.rf_ram.memory[129][2] ;
 wire \u_cpu.rf_ram.memory[129][3] ;
 wire \u_cpu.rf_ram.memory[129][4] ;
 wire \u_cpu.rf_ram.memory[129][5] ;
 wire \u_cpu.rf_ram.memory[129][6] ;
 wire \u_cpu.rf_ram.memory[129][7] ;
 wire \u_cpu.rf_ram.memory[12][0] ;
 wire \u_cpu.rf_ram.memory[12][1] ;
 wire \u_cpu.rf_ram.memory[12][2] ;
 wire \u_cpu.rf_ram.memory[12][3] ;
 wire \u_cpu.rf_ram.memory[12][4] ;
 wire \u_cpu.rf_ram.memory[12][5] ;
 wire \u_cpu.rf_ram.memory[12][6] ;
 wire \u_cpu.rf_ram.memory[12][7] ;
 wire \u_cpu.rf_ram.memory[130][0] ;
 wire \u_cpu.rf_ram.memory[130][1] ;
 wire \u_cpu.rf_ram.memory[130][2] ;
 wire \u_cpu.rf_ram.memory[130][3] ;
 wire \u_cpu.rf_ram.memory[130][4] ;
 wire \u_cpu.rf_ram.memory[130][5] ;
 wire \u_cpu.rf_ram.memory[130][6] ;
 wire \u_cpu.rf_ram.memory[130][7] ;
 wire \u_cpu.rf_ram.memory[131][0] ;
 wire \u_cpu.rf_ram.memory[131][1] ;
 wire \u_cpu.rf_ram.memory[131][2] ;
 wire \u_cpu.rf_ram.memory[131][3] ;
 wire \u_cpu.rf_ram.memory[131][4] ;
 wire \u_cpu.rf_ram.memory[131][5] ;
 wire \u_cpu.rf_ram.memory[131][6] ;
 wire \u_cpu.rf_ram.memory[131][7] ;
 wire \u_cpu.rf_ram.memory[132][0] ;
 wire \u_cpu.rf_ram.memory[132][1] ;
 wire \u_cpu.rf_ram.memory[132][2] ;
 wire \u_cpu.rf_ram.memory[132][3] ;
 wire \u_cpu.rf_ram.memory[132][4] ;
 wire \u_cpu.rf_ram.memory[132][5] ;
 wire \u_cpu.rf_ram.memory[132][6] ;
 wire \u_cpu.rf_ram.memory[132][7] ;
 wire \u_cpu.rf_ram.memory[133][0] ;
 wire \u_cpu.rf_ram.memory[133][1] ;
 wire \u_cpu.rf_ram.memory[133][2] ;
 wire \u_cpu.rf_ram.memory[133][3] ;
 wire \u_cpu.rf_ram.memory[133][4] ;
 wire \u_cpu.rf_ram.memory[133][5] ;
 wire \u_cpu.rf_ram.memory[133][6] ;
 wire \u_cpu.rf_ram.memory[133][7] ;
 wire \u_cpu.rf_ram.memory[134][0] ;
 wire \u_cpu.rf_ram.memory[134][1] ;
 wire \u_cpu.rf_ram.memory[134][2] ;
 wire \u_cpu.rf_ram.memory[134][3] ;
 wire \u_cpu.rf_ram.memory[134][4] ;
 wire \u_cpu.rf_ram.memory[134][5] ;
 wire \u_cpu.rf_ram.memory[134][6] ;
 wire \u_cpu.rf_ram.memory[134][7] ;
 wire \u_cpu.rf_ram.memory[135][0] ;
 wire \u_cpu.rf_ram.memory[135][1] ;
 wire \u_cpu.rf_ram.memory[135][2] ;
 wire \u_cpu.rf_ram.memory[135][3] ;
 wire \u_cpu.rf_ram.memory[135][4] ;
 wire \u_cpu.rf_ram.memory[135][5] ;
 wire \u_cpu.rf_ram.memory[135][6] ;
 wire \u_cpu.rf_ram.memory[135][7] ;
 wire \u_cpu.rf_ram.memory[136][0] ;
 wire \u_cpu.rf_ram.memory[136][1] ;
 wire \u_cpu.rf_ram.memory[136][2] ;
 wire \u_cpu.rf_ram.memory[136][3] ;
 wire \u_cpu.rf_ram.memory[136][4] ;
 wire \u_cpu.rf_ram.memory[136][5] ;
 wire \u_cpu.rf_ram.memory[136][6] ;
 wire \u_cpu.rf_ram.memory[136][7] ;
 wire \u_cpu.rf_ram.memory[137][0] ;
 wire \u_cpu.rf_ram.memory[137][1] ;
 wire \u_cpu.rf_ram.memory[137][2] ;
 wire \u_cpu.rf_ram.memory[137][3] ;
 wire \u_cpu.rf_ram.memory[137][4] ;
 wire \u_cpu.rf_ram.memory[137][5] ;
 wire \u_cpu.rf_ram.memory[137][6] ;
 wire \u_cpu.rf_ram.memory[137][7] ;
 wire \u_cpu.rf_ram.memory[138][0] ;
 wire \u_cpu.rf_ram.memory[138][1] ;
 wire \u_cpu.rf_ram.memory[138][2] ;
 wire \u_cpu.rf_ram.memory[138][3] ;
 wire \u_cpu.rf_ram.memory[138][4] ;
 wire \u_cpu.rf_ram.memory[138][5] ;
 wire \u_cpu.rf_ram.memory[138][6] ;
 wire \u_cpu.rf_ram.memory[138][7] ;
 wire \u_cpu.rf_ram.memory[139][0] ;
 wire \u_cpu.rf_ram.memory[139][1] ;
 wire \u_cpu.rf_ram.memory[139][2] ;
 wire \u_cpu.rf_ram.memory[139][3] ;
 wire \u_cpu.rf_ram.memory[139][4] ;
 wire \u_cpu.rf_ram.memory[139][5] ;
 wire \u_cpu.rf_ram.memory[139][6] ;
 wire \u_cpu.rf_ram.memory[139][7] ;
 wire \u_cpu.rf_ram.memory[13][0] ;
 wire \u_cpu.rf_ram.memory[13][1] ;
 wire \u_cpu.rf_ram.memory[13][2] ;
 wire \u_cpu.rf_ram.memory[13][3] ;
 wire \u_cpu.rf_ram.memory[13][4] ;
 wire \u_cpu.rf_ram.memory[13][5] ;
 wire \u_cpu.rf_ram.memory[13][6] ;
 wire \u_cpu.rf_ram.memory[13][7] ;
 wire \u_cpu.rf_ram.memory[140][0] ;
 wire \u_cpu.rf_ram.memory[140][1] ;
 wire \u_cpu.rf_ram.memory[140][2] ;
 wire \u_cpu.rf_ram.memory[140][3] ;
 wire \u_cpu.rf_ram.memory[140][4] ;
 wire \u_cpu.rf_ram.memory[140][5] ;
 wire \u_cpu.rf_ram.memory[140][6] ;
 wire \u_cpu.rf_ram.memory[140][7] ;
 wire \u_cpu.rf_ram.memory[141][0] ;
 wire \u_cpu.rf_ram.memory[141][1] ;
 wire \u_cpu.rf_ram.memory[141][2] ;
 wire \u_cpu.rf_ram.memory[141][3] ;
 wire \u_cpu.rf_ram.memory[141][4] ;
 wire \u_cpu.rf_ram.memory[141][5] ;
 wire \u_cpu.rf_ram.memory[141][6] ;
 wire \u_cpu.rf_ram.memory[141][7] ;
 wire \u_cpu.rf_ram.memory[142][0] ;
 wire \u_cpu.rf_ram.memory[142][1] ;
 wire \u_cpu.rf_ram.memory[142][2] ;
 wire \u_cpu.rf_ram.memory[142][3] ;
 wire \u_cpu.rf_ram.memory[142][4] ;
 wire \u_cpu.rf_ram.memory[142][5] ;
 wire \u_cpu.rf_ram.memory[142][6] ;
 wire \u_cpu.rf_ram.memory[142][7] ;
 wire \u_cpu.rf_ram.memory[143][0] ;
 wire \u_cpu.rf_ram.memory[143][1] ;
 wire \u_cpu.rf_ram.memory[143][2] ;
 wire \u_cpu.rf_ram.memory[143][3] ;
 wire \u_cpu.rf_ram.memory[143][4] ;
 wire \u_cpu.rf_ram.memory[143][5] ;
 wire \u_cpu.rf_ram.memory[143][6] ;
 wire \u_cpu.rf_ram.memory[143][7] ;
 wire \u_cpu.rf_ram.memory[14][0] ;
 wire \u_cpu.rf_ram.memory[14][1] ;
 wire \u_cpu.rf_ram.memory[14][2] ;
 wire \u_cpu.rf_ram.memory[14][3] ;
 wire \u_cpu.rf_ram.memory[14][4] ;
 wire \u_cpu.rf_ram.memory[14][5] ;
 wire \u_cpu.rf_ram.memory[14][6] ;
 wire \u_cpu.rf_ram.memory[14][7] ;
 wire \u_cpu.rf_ram.memory[15][0] ;
 wire \u_cpu.rf_ram.memory[15][1] ;
 wire \u_cpu.rf_ram.memory[15][2] ;
 wire \u_cpu.rf_ram.memory[15][3] ;
 wire \u_cpu.rf_ram.memory[15][4] ;
 wire \u_cpu.rf_ram.memory[15][5] ;
 wire \u_cpu.rf_ram.memory[15][6] ;
 wire \u_cpu.rf_ram.memory[15][7] ;
 wire \u_cpu.rf_ram.memory[16][0] ;
 wire \u_cpu.rf_ram.memory[16][1] ;
 wire \u_cpu.rf_ram.memory[16][2] ;
 wire \u_cpu.rf_ram.memory[16][3] ;
 wire \u_cpu.rf_ram.memory[16][4] ;
 wire \u_cpu.rf_ram.memory[16][5] ;
 wire \u_cpu.rf_ram.memory[16][6] ;
 wire \u_cpu.rf_ram.memory[16][7] ;
 wire \u_cpu.rf_ram.memory[17][0] ;
 wire \u_cpu.rf_ram.memory[17][1] ;
 wire \u_cpu.rf_ram.memory[17][2] ;
 wire \u_cpu.rf_ram.memory[17][3] ;
 wire \u_cpu.rf_ram.memory[17][4] ;
 wire \u_cpu.rf_ram.memory[17][5] ;
 wire \u_cpu.rf_ram.memory[17][6] ;
 wire \u_cpu.rf_ram.memory[17][7] ;
 wire \u_cpu.rf_ram.memory[18][0] ;
 wire \u_cpu.rf_ram.memory[18][1] ;
 wire \u_cpu.rf_ram.memory[18][2] ;
 wire \u_cpu.rf_ram.memory[18][3] ;
 wire \u_cpu.rf_ram.memory[18][4] ;
 wire \u_cpu.rf_ram.memory[18][5] ;
 wire \u_cpu.rf_ram.memory[18][6] ;
 wire \u_cpu.rf_ram.memory[18][7] ;
 wire \u_cpu.rf_ram.memory[19][0] ;
 wire \u_cpu.rf_ram.memory[19][1] ;
 wire \u_cpu.rf_ram.memory[19][2] ;
 wire \u_cpu.rf_ram.memory[19][3] ;
 wire \u_cpu.rf_ram.memory[19][4] ;
 wire \u_cpu.rf_ram.memory[19][5] ;
 wire \u_cpu.rf_ram.memory[19][6] ;
 wire \u_cpu.rf_ram.memory[19][7] ;
 wire \u_cpu.rf_ram.memory[1][0] ;
 wire \u_cpu.rf_ram.memory[1][1] ;
 wire \u_cpu.rf_ram.memory[1][2] ;
 wire \u_cpu.rf_ram.memory[1][3] ;
 wire \u_cpu.rf_ram.memory[1][4] ;
 wire \u_cpu.rf_ram.memory[1][5] ;
 wire \u_cpu.rf_ram.memory[1][6] ;
 wire \u_cpu.rf_ram.memory[1][7] ;
 wire \u_cpu.rf_ram.memory[20][0] ;
 wire \u_cpu.rf_ram.memory[20][1] ;
 wire \u_cpu.rf_ram.memory[20][2] ;
 wire \u_cpu.rf_ram.memory[20][3] ;
 wire \u_cpu.rf_ram.memory[20][4] ;
 wire \u_cpu.rf_ram.memory[20][5] ;
 wire \u_cpu.rf_ram.memory[20][6] ;
 wire \u_cpu.rf_ram.memory[20][7] ;
 wire \u_cpu.rf_ram.memory[21][0] ;
 wire \u_cpu.rf_ram.memory[21][1] ;
 wire \u_cpu.rf_ram.memory[21][2] ;
 wire \u_cpu.rf_ram.memory[21][3] ;
 wire \u_cpu.rf_ram.memory[21][4] ;
 wire \u_cpu.rf_ram.memory[21][5] ;
 wire \u_cpu.rf_ram.memory[21][6] ;
 wire \u_cpu.rf_ram.memory[21][7] ;
 wire \u_cpu.rf_ram.memory[22][0] ;
 wire \u_cpu.rf_ram.memory[22][1] ;
 wire \u_cpu.rf_ram.memory[22][2] ;
 wire \u_cpu.rf_ram.memory[22][3] ;
 wire \u_cpu.rf_ram.memory[22][4] ;
 wire \u_cpu.rf_ram.memory[22][5] ;
 wire \u_cpu.rf_ram.memory[22][6] ;
 wire \u_cpu.rf_ram.memory[22][7] ;
 wire \u_cpu.rf_ram.memory[23][0] ;
 wire \u_cpu.rf_ram.memory[23][1] ;
 wire \u_cpu.rf_ram.memory[23][2] ;
 wire \u_cpu.rf_ram.memory[23][3] ;
 wire \u_cpu.rf_ram.memory[23][4] ;
 wire \u_cpu.rf_ram.memory[23][5] ;
 wire \u_cpu.rf_ram.memory[23][6] ;
 wire \u_cpu.rf_ram.memory[23][7] ;
 wire \u_cpu.rf_ram.memory[24][0] ;
 wire \u_cpu.rf_ram.memory[24][1] ;
 wire \u_cpu.rf_ram.memory[24][2] ;
 wire \u_cpu.rf_ram.memory[24][3] ;
 wire \u_cpu.rf_ram.memory[24][4] ;
 wire \u_cpu.rf_ram.memory[24][5] ;
 wire \u_cpu.rf_ram.memory[24][6] ;
 wire \u_cpu.rf_ram.memory[24][7] ;
 wire \u_cpu.rf_ram.memory[25][0] ;
 wire \u_cpu.rf_ram.memory[25][1] ;
 wire \u_cpu.rf_ram.memory[25][2] ;
 wire \u_cpu.rf_ram.memory[25][3] ;
 wire \u_cpu.rf_ram.memory[25][4] ;
 wire \u_cpu.rf_ram.memory[25][5] ;
 wire \u_cpu.rf_ram.memory[25][6] ;
 wire \u_cpu.rf_ram.memory[25][7] ;
 wire \u_cpu.rf_ram.memory[26][0] ;
 wire \u_cpu.rf_ram.memory[26][1] ;
 wire \u_cpu.rf_ram.memory[26][2] ;
 wire \u_cpu.rf_ram.memory[26][3] ;
 wire \u_cpu.rf_ram.memory[26][4] ;
 wire \u_cpu.rf_ram.memory[26][5] ;
 wire \u_cpu.rf_ram.memory[26][6] ;
 wire \u_cpu.rf_ram.memory[26][7] ;
 wire \u_cpu.rf_ram.memory[27][0] ;
 wire \u_cpu.rf_ram.memory[27][1] ;
 wire \u_cpu.rf_ram.memory[27][2] ;
 wire \u_cpu.rf_ram.memory[27][3] ;
 wire \u_cpu.rf_ram.memory[27][4] ;
 wire \u_cpu.rf_ram.memory[27][5] ;
 wire \u_cpu.rf_ram.memory[27][6] ;
 wire \u_cpu.rf_ram.memory[27][7] ;
 wire \u_cpu.rf_ram.memory[28][0] ;
 wire \u_cpu.rf_ram.memory[28][1] ;
 wire \u_cpu.rf_ram.memory[28][2] ;
 wire \u_cpu.rf_ram.memory[28][3] ;
 wire \u_cpu.rf_ram.memory[28][4] ;
 wire \u_cpu.rf_ram.memory[28][5] ;
 wire \u_cpu.rf_ram.memory[28][6] ;
 wire \u_cpu.rf_ram.memory[28][7] ;
 wire \u_cpu.rf_ram.memory[29][0] ;
 wire \u_cpu.rf_ram.memory[29][1] ;
 wire \u_cpu.rf_ram.memory[29][2] ;
 wire \u_cpu.rf_ram.memory[29][3] ;
 wire \u_cpu.rf_ram.memory[29][4] ;
 wire \u_cpu.rf_ram.memory[29][5] ;
 wire \u_cpu.rf_ram.memory[29][6] ;
 wire \u_cpu.rf_ram.memory[29][7] ;
 wire \u_cpu.rf_ram.memory[2][0] ;
 wire \u_cpu.rf_ram.memory[2][1] ;
 wire \u_cpu.rf_ram.memory[2][2] ;
 wire \u_cpu.rf_ram.memory[2][3] ;
 wire \u_cpu.rf_ram.memory[2][4] ;
 wire \u_cpu.rf_ram.memory[2][5] ;
 wire \u_cpu.rf_ram.memory[2][6] ;
 wire \u_cpu.rf_ram.memory[2][7] ;
 wire \u_cpu.rf_ram.memory[30][0] ;
 wire \u_cpu.rf_ram.memory[30][1] ;
 wire \u_cpu.rf_ram.memory[30][2] ;
 wire \u_cpu.rf_ram.memory[30][3] ;
 wire \u_cpu.rf_ram.memory[30][4] ;
 wire \u_cpu.rf_ram.memory[30][5] ;
 wire \u_cpu.rf_ram.memory[30][6] ;
 wire \u_cpu.rf_ram.memory[30][7] ;
 wire \u_cpu.rf_ram.memory[31][0] ;
 wire \u_cpu.rf_ram.memory[31][1] ;
 wire \u_cpu.rf_ram.memory[31][2] ;
 wire \u_cpu.rf_ram.memory[31][3] ;
 wire \u_cpu.rf_ram.memory[31][4] ;
 wire \u_cpu.rf_ram.memory[31][5] ;
 wire \u_cpu.rf_ram.memory[31][6] ;
 wire \u_cpu.rf_ram.memory[31][7] ;
 wire \u_cpu.rf_ram.memory[32][0] ;
 wire \u_cpu.rf_ram.memory[32][1] ;
 wire \u_cpu.rf_ram.memory[32][2] ;
 wire \u_cpu.rf_ram.memory[32][3] ;
 wire \u_cpu.rf_ram.memory[32][4] ;
 wire \u_cpu.rf_ram.memory[32][5] ;
 wire \u_cpu.rf_ram.memory[32][6] ;
 wire \u_cpu.rf_ram.memory[32][7] ;
 wire \u_cpu.rf_ram.memory[33][0] ;
 wire \u_cpu.rf_ram.memory[33][1] ;
 wire \u_cpu.rf_ram.memory[33][2] ;
 wire \u_cpu.rf_ram.memory[33][3] ;
 wire \u_cpu.rf_ram.memory[33][4] ;
 wire \u_cpu.rf_ram.memory[33][5] ;
 wire \u_cpu.rf_ram.memory[33][6] ;
 wire \u_cpu.rf_ram.memory[33][7] ;
 wire \u_cpu.rf_ram.memory[34][0] ;
 wire \u_cpu.rf_ram.memory[34][1] ;
 wire \u_cpu.rf_ram.memory[34][2] ;
 wire \u_cpu.rf_ram.memory[34][3] ;
 wire \u_cpu.rf_ram.memory[34][4] ;
 wire \u_cpu.rf_ram.memory[34][5] ;
 wire \u_cpu.rf_ram.memory[34][6] ;
 wire \u_cpu.rf_ram.memory[34][7] ;
 wire \u_cpu.rf_ram.memory[35][0] ;
 wire \u_cpu.rf_ram.memory[35][1] ;
 wire \u_cpu.rf_ram.memory[35][2] ;
 wire \u_cpu.rf_ram.memory[35][3] ;
 wire \u_cpu.rf_ram.memory[35][4] ;
 wire \u_cpu.rf_ram.memory[35][5] ;
 wire \u_cpu.rf_ram.memory[35][6] ;
 wire \u_cpu.rf_ram.memory[35][7] ;
 wire \u_cpu.rf_ram.memory[36][0] ;
 wire \u_cpu.rf_ram.memory[36][1] ;
 wire \u_cpu.rf_ram.memory[36][2] ;
 wire \u_cpu.rf_ram.memory[36][3] ;
 wire \u_cpu.rf_ram.memory[36][4] ;
 wire \u_cpu.rf_ram.memory[36][5] ;
 wire \u_cpu.rf_ram.memory[36][6] ;
 wire \u_cpu.rf_ram.memory[36][7] ;
 wire \u_cpu.rf_ram.memory[37][0] ;
 wire \u_cpu.rf_ram.memory[37][1] ;
 wire \u_cpu.rf_ram.memory[37][2] ;
 wire \u_cpu.rf_ram.memory[37][3] ;
 wire \u_cpu.rf_ram.memory[37][4] ;
 wire \u_cpu.rf_ram.memory[37][5] ;
 wire \u_cpu.rf_ram.memory[37][6] ;
 wire \u_cpu.rf_ram.memory[37][7] ;
 wire \u_cpu.rf_ram.memory[38][0] ;
 wire \u_cpu.rf_ram.memory[38][1] ;
 wire \u_cpu.rf_ram.memory[38][2] ;
 wire \u_cpu.rf_ram.memory[38][3] ;
 wire \u_cpu.rf_ram.memory[38][4] ;
 wire \u_cpu.rf_ram.memory[38][5] ;
 wire \u_cpu.rf_ram.memory[38][6] ;
 wire \u_cpu.rf_ram.memory[38][7] ;
 wire \u_cpu.rf_ram.memory[39][0] ;
 wire \u_cpu.rf_ram.memory[39][1] ;
 wire \u_cpu.rf_ram.memory[39][2] ;
 wire \u_cpu.rf_ram.memory[39][3] ;
 wire \u_cpu.rf_ram.memory[39][4] ;
 wire \u_cpu.rf_ram.memory[39][5] ;
 wire \u_cpu.rf_ram.memory[39][6] ;
 wire \u_cpu.rf_ram.memory[39][7] ;
 wire \u_cpu.rf_ram.memory[3][0] ;
 wire \u_cpu.rf_ram.memory[3][1] ;
 wire \u_cpu.rf_ram.memory[3][2] ;
 wire \u_cpu.rf_ram.memory[3][3] ;
 wire \u_cpu.rf_ram.memory[3][4] ;
 wire \u_cpu.rf_ram.memory[3][5] ;
 wire \u_cpu.rf_ram.memory[3][6] ;
 wire \u_cpu.rf_ram.memory[3][7] ;
 wire \u_cpu.rf_ram.memory[40][0] ;
 wire \u_cpu.rf_ram.memory[40][1] ;
 wire \u_cpu.rf_ram.memory[40][2] ;
 wire \u_cpu.rf_ram.memory[40][3] ;
 wire \u_cpu.rf_ram.memory[40][4] ;
 wire \u_cpu.rf_ram.memory[40][5] ;
 wire \u_cpu.rf_ram.memory[40][6] ;
 wire \u_cpu.rf_ram.memory[40][7] ;
 wire \u_cpu.rf_ram.memory[41][0] ;
 wire \u_cpu.rf_ram.memory[41][1] ;
 wire \u_cpu.rf_ram.memory[41][2] ;
 wire \u_cpu.rf_ram.memory[41][3] ;
 wire \u_cpu.rf_ram.memory[41][4] ;
 wire \u_cpu.rf_ram.memory[41][5] ;
 wire \u_cpu.rf_ram.memory[41][6] ;
 wire \u_cpu.rf_ram.memory[41][7] ;
 wire \u_cpu.rf_ram.memory[42][0] ;
 wire \u_cpu.rf_ram.memory[42][1] ;
 wire \u_cpu.rf_ram.memory[42][2] ;
 wire \u_cpu.rf_ram.memory[42][3] ;
 wire \u_cpu.rf_ram.memory[42][4] ;
 wire \u_cpu.rf_ram.memory[42][5] ;
 wire \u_cpu.rf_ram.memory[42][6] ;
 wire \u_cpu.rf_ram.memory[42][7] ;
 wire \u_cpu.rf_ram.memory[43][0] ;
 wire \u_cpu.rf_ram.memory[43][1] ;
 wire \u_cpu.rf_ram.memory[43][2] ;
 wire \u_cpu.rf_ram.memory[43][3] ;
 wire \u_cpu.rf_ram.memory[43][4] ;
 wire \u_cpu.rf_ram.memory[43][5] ;
 wire \u_cpu.rf_ram.memory[43][6] ;
 wire \u_cpu.rf_ram.memory[43][7] ;
 wire \u_cpu.rf_ram.memory[44][0] ;
 wire \u_cpu.rf_ram.memory[44][1] ;
 wire \u_cpu.rf_ram.memory[44][2] ;
 wire \u_cpu.rf_ram.memory[44][3] ;
 wire \u_cpu.rf_ram.memory[44][4] ;
 wire \u_cpu.rf_ram.memory[44][5] ;
 wire \u_cpu.rf_ram.memory[44][6] ;
 wire \u_cpu.rf_ram.memory[44][7] ;
 wire \u_cpu.rf_ram.memory[45][0] ;
 wire \u_cpu.rf_ram.memory[45][1] ;
 wire \u_cpu.rf_ram.memory[45][2] ;
 wire \u_cpu.rf_ram.memory[45][3] ;
 wire \u_cpu.rf_ram.memory[45][4] ;
 wire \u_cpu.rf_ram.memory[45][5] ;
 wire \u_cpu.rf_ram.memory[45][6] ;
 wire \u_cpu.rf_ram.memory[45][7] ;
 wire \u_cpu.rf_ram.memory[46][0] ;
 wire \u_cpu.rf_ram.memory[46][1] ;
 wire \u_cpu.rf_ram.memory[46][2] ;
 wire \u_cpu.rf_ram.memory[46][3] ;
 wire \u_cpu.rf_ram.memory[46][4] ;
 wire \u_cpu.rf_ram.memory[46][5] ;
 wire \u_cpu.rf_ram.memory[46][6] ;
 wire \u_cpu.rf_ram.memory[46][7] ;
 wire \u_cpu.rf_ram.memory[47][0] ;
 wire \u_cpu.rf_ram.memory[47][1] ;
 wire \u_cpu.rf_ram.memory[47][2] ;
 wire \u_cpu.rf_ram.memory[47][3] ;
 wire \u_cpu.rf_ram.memory[47][4] ;
 wire \u_cpu.rf_ram.memory[47][5] ;
 wire \u_cpu.rf_ram.memory[47][6] ;
 wire \u_cpu.rf_ram.memory[47][7] ;
 wire \u_cpu.rf_ram.memory[48][0] ;
 wire \u_cpu.rf_ram.memory[48][1] ;
 wire \u_cpu.rf_ram.memory[48][2] ;
 wire \u_cpu.rf_ram.memory[48][3] ;
 wire \u_cpu.rf_ram.memory[48][4] ;
 wire \u_cpu.rf_ram.memory[48][5] ;
 wire \u_cpu.rf_ram.memory[48][6] ;
 wire \u_cpu.rf_ram.memory[48][7] ;
 wire \u_cpu.rf_ram.memory[49][0] ;
 wire \u_cpu.rf_ram.memory[49][1] ;
 wire \u_cpu.rf_ram.memory[49][2] ;
 wire \u_cpu.rf_ram.memory[49][3] ;
 wire \u_cpu.rf_ram.memory[49][4] ;
 wire \u_cpu.rf_ram.memory[49][5] ;
 wire \u_cpu.rf_ram.memory[49][6] ;
 wire \u_cpu.rf_ram.memory[49][7] ;
 wire \u_cpu.rf_ram.memory[4][0] ;
 wire \u_cpu.rf_ram.memory[4][1] ;
 wire \u_cpu.rf_ram.memory[4][2] ;
 wire \u_cpu.rf_ram.memory[4][3] ;
 wire \u_cpu.rf_ram.memory[4][4] ;
 wire \u_cpu.rf_ram.memory[4][5] ;
 wire \u_cpu.rf_ram.memory[4][6] ;
 wire \u_cpu.rf_ram.memory[4][7] ;
 wire \u_cpu.rf_ram.memory[50][0] ;
 wire \u_cpu.rf_ram.memory[50][1] ;
 wire \u_cpu.rf_ram.memory[50][2] ;
 wire \u_cpu.rf_ram.memory[50][3] ;
 wire \u_cpu.rf_ram.memory[50][4] ;
 wire \u_cpu.rf_ram.memory[50][5] ;
 wire \u_cpu.rf_ram.memory[50][6] ;
 wire \u_cpu.rf_ram.memory[50][7] ;
 wire \u_cpu.rf_ram.memory[51][0] ;
 wire \u_cpu.rf_ram.memory[51][1] ;
 wire \u_cpu.rf_ram.memory[51][2] ;
 wire \u_cpu.rf_ram.memory[51][3] ;
 wire \u_cpu.rf_ram.memory[51][4] ;
 wire \u_cpu.rf_ram.memory[51][5] ;
 wire \u_cpu.rf_ram.memory[51][6] ;
 wire \u_cpu.rf_ram.memory[51][7] ;
 wire \u_cpu.rf_ram.memory[52][0] ;
 wire \u_cpu.rf_ram.memory[52][1] ;
 wire \u_cpu.rf_ram.memory[52][2] ;
 wire \u_cpu.rf_ram.memory[52][3] ;
 wire \u_cpu.rf_ram.memory[52][4] ;
 wire \u_cpu.rf_ram.memory[52][5] ;
 wire \u_cpu.rf_ram.memory[52][6] ;
 wire \u_cpu.rf_ram.memory[52][7] ;
 wire \u_cpu.rf_ram.memory[53][0] ;
 wire \u_cpu.rf_ram.memory[53][1] ;
 wire \u_cpu.rf_ram.memory[53][2] ;
 wire \u_cpu.rf_ram.memory[53][3] ;
 wire \u_cpu.rf_ram.memory[53][4] ;
 wire \u_cpu.rf_ram.memory[53][5] ;
 wire \u_cpu.rf_ram.memory[53][6] ;
 wire \u_cpu.rf_ram.memory[53][7] ;
 wire \u_cpu.rf_ram.memory[54][0] ;
 wire \u_cpu.rf_ram.memory[54][1] ;
 wire \u_cpu.rf_ram.memory[54][2] ;
 wire \u_cpu.rf_ram.memory[54][3] ;
 wire \u_cpu.rf_ram.memory[54][4] ;
 wire \u_cpu.rf_ram.memory[54][5] ;
 wire \u_cpu.rf_ram.memory[54][6] ;
 wire \u_cpu.rf_ram.memory[54][7] ;
 wire \u_cpu.rf_ram.memory[55][0] ;
 wire \u_cpu.rf_ram.memory[55][1] ;
 wire \u_cpu.rf_ram.memory[55][2] ;
 wire \u_cpu.rf_ram.memory[55][3] ;
 wire \u_cpu.rf_ram.memory[55][4] ;
 wire \u_cpu.rf_ram.memory[55][5] ;
 wire \u_cpu.rf_ram.memory[55][6] ;
 wire \u_cpu.rf_ram.memory[55][7] ;
 wire \u_cpu.rf_ram.memory[56][0] ;
 wire \u_cpu.rf_ram.memory[56][1] ;
 wire \u_cpu.rf_ram.memory[56][2] ;
 wire \u_cpu.rf_ram.memory[56][3] ;
 wire \u_cpu.rf_ram.memory[56][4] ;
 wire \u_cpu.rf_ram.memory[56][5] ;
 wire \u_cpu.rf_ram.memory[56][6] ;
 wire \u_cpu.rf_ram.memory[56][7] ;
 wire \u_cpu.rf_ram.memory[57][0] ;
 wire \u_cpu.rf_ram.memory[57][1] ;
 wire \u_cpu.rf_ram.memory[57][2] ;
 wire \u_cpu.rf_ram.memory[57][3] ;
 wire \u_cpu.rf_ram.memory[57][4] ;
 wire \u_cpu.rf_ram.memory[57][5] ;
 wire \u_cpu.rf_ram.memory[57][6] ;
 wire \u_cpu.rf_ram.memory[57][7] ;
 wire \u_cpu.rf_ram.memory[58][0] ;
 wire \u_cpu.rf_ram.memory[58][1] ;
 wire \u_cpu.rf_ram.memory[58][2] ;
 wire \u_cpu.rf_ram.memory[58][3] ;
 wire \u_cpu.rf_ram.memory[58][4] ;
 wire \u_cpu.rf_ram.memory[58][5] ;
 wire \u_cpu.rf_ram.memory[58][6] ;
 wire \u_cpu.rf_ram.memory[58][7] ;
 wire \u_cpu.rf_ram.memory[59][0] ;
 wire \u_cpu.rf_ram.memory[59][1] ;
 wire \u_cpu.rf_ram.memory[59][2] ;
 wire \u_cpu.rf_ram.memory[59][3] ;
 wire \u_cpu.rf_ram.memory[59][4] ;
 wire \u_cpu.rf_ram.memory[59][5] ;
 wire \u_cpu.rf_ram.memory[59][6] ;
 wire \u_cpu.rf_ram.memory[59][7] ;
 wire \u_cpu.rf_ram.memory[5][0] ;
 wire \u_cpu.rf_ram.memory[5][1] ;
 wire \u_cpu.rf_ram.memory[5][2] ;
 wire \u_cpu.rf_ram.memory[5][3] ;
 wire \u_cpu.rf_ram.memory[5][4] ;
 wire \u_cpu.rf_ram.memory[5][5] ;
 wire \u_cpu.rf_ram.memory[5][6] ;
 wire \u_cpu.rf_ram.memory[5][7] ;
 wire \u_cpu.rf_ram.memory[60][0] ;
 wire \u_cpu.rf_ram.memory[60][1] ;
 wire \u_cpu.rf_ram.memory[60][2] ;
 wire \u_cpu.rf_ram.memory[60][3] ;
 wire \u_cpu.rf_ram.memory[60][4] ;
 wire \u_cpu.rf_ram.memory[60][5] ;
 wire \u_cpu.rf_ram.memory[60][6] ;
 wire \u_cpu.rf_ram.memory[60][7] ;
 wire \u_cpu.rf_ram.memory[61][0] ;
 wire \u_cpu.rf_ram.memory[61][1] ;
 wire \u_cpu.rf_ram.memory[61][2] ;
 wire \u_cpu.rf_ram.memory[61][3] ;
 wire \u_cpu.rf_ram.memory[61][4] ;
 wire \u_cpu.rf_ram.memory[61][5] ;
 wire \u_cpu.rf_ram.memory[61][6] ;
 wire \u_cpu.rf_ram.memory[61][7] ;
 wire \u_cpu.rf_ram.memory[62][0] ;
 wire \u_cpu.rf_ram.memory[62][1] ;
 wire \u_cpu.rf_ram.memory[62][2] ;
 wire \u_cpu.rf_ram.memory[62][3] ;
 wire \u_cpu.rf_ram.memory[62][4] ;
 wire \u_cpu.rf_ram.memory[62][5] ;
 wire \u_cpu.rf_ram.memory[62][6] ;
 wire \u_cpu.rf_ram.memory[62][7] ;
 wire \u_cpu.rf_ram.memory[63][0] ;
 wire \u_cpu.rf_ram.memory[63][1] ;
 wire \u_cpu.rf_ram.memory[63][2] ;
 wire \u_cpu.rf_ram.memory[63][3] ;
 wire \u_cpu.rf_ram.memory[63][4] ;
 wire \u_cpu.rf_ram.memory[63][5] ;
 wire \u_cpu.rf_ram.memory[63][6] ;
 wire \u_cpu.rf_ram.memory[63][7] ;
 wire \u_cpu.rf_ram.memory[64][0] ;
 wire \u_cpu.rf_ram.memory[64][1] ;
 wire \u_cpu.rf_ram.memory[64][2] ;
 wire \u_cpu.rf_ram.memory[64][3] ;
 wire \u_cpu.rf_ram.memory[64][4] ;
 wire \u_cpu.rf_ram.memory[64][5] ;
 wire \u_cpu.rf_ram.memory[64][6] ;
 wire \u_cpu.rf_ram.memory[64][7] ;
 wire \u_cpu.rf_ram.memory[65][0] ;
 wire \u_cpu.rf_ram.memory[65][1] ;
 wire \u_cpu.rf_ram.memory[65][2] ;
 wire \u_cpu.rf_ram.memory[65][3] ;
 wire \u_cpu.rf_ram.memory[65][4] ;
 wire \u_cpu.rf_ram.memory[65][5] ;
 wire \u_cpu.rf_ram.memory[65][6] ;
 wire \u_cpu.rf_ram.memory[65][7] ;
 wire \u_cpu.rf_ram.memory[66][0] ;
 wire \u_cpu.rf_ram.memory[66][1] ;
 wire \u_cpu.rf_ram.memory[66][2] ;
 wire \u_cpu.rf_ram.memory[66][3] ;
 wire \u_cpu.rf_ram.memory[66][4] ;
 wire \u_cpu.rf_ram.memory[66][5] ;
 wire \u_cpu.rf_ram.memory[66][6] ;
 wire \u_cpu.rf_ram.memory[66][7] ;
 wire \u_cpu.rf_ram.memory[67][0] ;
 wire \u_cpu.rf_ram.memory[67][1] ;
 wire \u_cpu.rf_ram.memory[67][2] ;
 wire \u_cpu.rf_ram.memory[67][3] ;
 wire \u_cpu.rf_ram.memory[67][4] ;
 wire \u_cpu.rf_ram.memory[67][5] ;
 wire \u_cpu.rf_ram.memory[67][6] ;
 wire \u_cpu.rf_ram.memory[67][7] ;
 wire \u_cpu.rf_ram.memory[68][0] ;
 wire \u_cpu.rf_ram.memory[68][1] ;
 wire \u_cpu.rf_ram.memory[68][2] ;
 wire \u_cpu.rf_ram.memory[68][3] ;
 wire \u_cpu.rf_ram.memory[68][4] ;
 wire \u_cpu.rf_ram.memory[68][5] ;
 wire \u_cpu.rf_ram.memory[68][6] ;
 wire \u_cpu.rf_ram.memory[68][7] ;
 wire \u_cpu.rf_ram.memory[69][0] ;
 wire \u_cpu.rf_ram.memory[69][1] ;
 wire \u_cpu.rf_ram.memory[69][2] ;
 wire \u_cpu.rf_ram.memory[69][3] ;
 wire \u_cpu.rf_ram.memory[69][4] ;
 wire \u_cpu.rf_ram.memory[69][5] ;
 wire \u_cpu.rf_ram.memory[69][6] ;
 wire \u_cpu.rf_ram.memory[69][7] ;
 wire \u_cpu.rf_ram.memory[6][0] ;
 wire \u_cpu.rf_ram.memory[6][1] ;
 wire \u_cpu.rf_ram.memory[6][2] ;
 wire \u_cpu.rf_ram.memory[6][3] ;
 wire \u_cpu.rf_ram.memory[6][4] ;
 wire \u_cpu.rf_ram.memory[6][5] ;
 wire \u_cpu.rf_ram.memory[6][6] ;
 wire \u_cpu.rf_ram.memory[6][7] ;
 wire \u_cpu.rf_ram.memory[70][0] ;
 wire \u_cpu.rf_ram.memory[70][1] ;
 wire \u_cpu.rf_ram.memory[70][2] ;
 wire \u_cpu.rf_ram.memory[70][3] ;
 wire \u_cpu.rf_ram.memory[70][4] ;
 wire \u_cpu.rf_ram.memory[70][5] ;
 wire \u_cpu.rf_ram.memory[70][6] ;
 wire \u_cpu.rf_ram.memory[70][7] ;
 wire \u_cpu.rf_ram.memory[71][0] ;
 wire \u_cpu.rf_ram.memory[71][1] ;
 wire \u_cpu.rf_ram.memory[71][2] ;
 wire \u_cpu.rf_ram.memory[71][3] ;
 wire \u_cpu.rf_ram.memory[71][4] ;
 wire \u_cpu.rf_ram.memory[71][5] ;
 wire \u_cpu.rf_ram.memory[71][6] ;
 wire \u_cpu.rf_ram.memory[71][7] ;
 wire \u_cpu.rf_ram.memory[72][0] ;
 wire \u_cpu.rf_ram.memory[72][1] ;
 wire \u_cpu.rf_ram.memory[72][2] ;
 wire \u_cpu.rf_ram.memory[72][3] ;
 wire \u_cpu.rf_ram.memory[72][4] ;
 wire \u_cpu.rf_ram.memory[72][5] ;
 wire \u_cpu.rf_ram.memory[72][6] ;
 wire \u_cpu.rf_ram.memory[72][7] ;
 wire \u_cpu.rf_ram.memory[73][0] ;
 wire \u_cpu.rf_ram.memory[73][1] ;
 wire \u_cpu.rf_ram.memory[73][2] ;
 wire \u_cpu.rf_ram.memory[73][3] ;
 wire \u_cpu.rf_ram.memory[73][4] ;
 wire \u_cpu.rf_ram.memory[73][5] ;
 wire \u_cpu.rf_ram.memory[73][6] ;
 wire \u_cpu.rf_ram.memory[73][7] ;
 wire \u_cpu.rf_ram.memory[74][0] ;
 wire \u_cpu.rf_ram.memory[74][1] ;
 wire \u_cpu.rf_ram.memory[74][2] ;
 wire \u_cpu.rf_ram.memory[74][3] ;
 wire \u_cpu.rf_ram.memory[74][4] ;
 wire \u_cpu.rf_ram.memory[74][5] ;
 wire \u_cpu.rf_ram.memory[74][6] ;
 wire \u_cpu.rf_ram.memory[74][7] ;
 wire \u_cpu.rf_ram.memory[75][0] ;
 wire \u_cpu.rf_ram.memory[75][1] ;
 wire \u_cpu.rf_ram.memory[75][2] ;
 wire \u_cpu.rf_ram.memory[75][3] ;
 wire \u_cpu.rf_ram.memory[75][4] ;
 wire \u_cpu.rf_ram.memory[75][5] ;
 wire \u_cpu.rf_ram.memory[75][6] ;
 wire \u_cpu.rf_ram.memory[75][7] ;
 wire \u_cpu.rf_ram.memory[76][0] ;
 wire \u_cpu.rf_ram.memory[76][1] ;
 wire \u_cpu.rf_ram.memory[76][2] ;
 wire \u_cpu.rf_ram.memory[76][3] ;
 wire \u_cpu.rf_ram.memory[76][4] ;
 wire \u_cpu.rf_ram.memory[76][5] ;
 wire \u_cpu.rf_ram.memory[76][6] ;
 wire \u_cpu.rf_ram.memory[76][7] ;
 wire \u_cpu.rf_ram.memory[77][0] ;
 wire \u_cpu.rf_ram.memory[77][1] ;
 wire \u_cpu.rf_ram.memory[77][2] ;
 wire \u_cpu.rf_ram.memory[77][3] ;
 wire \u_cpu.rf_ram.memory[77][4] ;
 wire \u_cpu.rf_ram.memory[77][5] ;
 wire \u_cpu.rf_ram.memory[77][6] ;
 wire \u_cpu.rf_ram.memory[77][7] ;
 wire \u_cpu.rf_ram.memory[78][0] ;
 wire \u_cpu.rf_ram.memory[78][1] ;
 wire \u_cpu.rf_ram.memory[78][2] ;
 wire \u_cpu.rf_ram.memory[78][3] ;
 wire \u_cpu.rf_ram.memory[78][4] ;
 wire \u_cpu.rf_ram.memory[78][5] ;
 wire \u_cpu.rf_ram.memory[78][6] ;
 wire \u_cpu.rf_ram.memory[78][7] ;
 wire \u_cpu.rf_ram.memory[79][0] ;
 wire \u_cpu.rf_ram.memory[79][1] ;
 wire \u_cpu.rf_ram.memory[79][2] ;
 wire \u_cpu.rf_ram.memory[79][3] ;
 wire \u_cpu.rf_ram.memory[79][4] ;
 wire \u_cpu.rf_ram.memory[79][5] ;
 wire \u_cpu.rf_ram.memory[79][6] ;
 wire \u_cpu.rf_ram.memory[79][7] ;
 wire \u_cpu.rf_ram.memory[7][0] ;
 wire \u_cpu.rf_ram.memory[7][1] ;
 wire \u_cpu.rf_ram.memory[7][2] ;
 wire \u_cpu.rf_ram.memory[7][3] ;
 wire \u_cpu.rf_ram.memory[7][4] ;
 wire \u_cpu.rf_ram.memory[7][5] ;
 wire \u_cpu.rf_ram.memory[7][6] ;
 wire \u_cpu.rf_ram.memory[7][7] ;
 wire \u_cpu.rf_ram.memory[80][0] ;
 wire \u_cpu.rf_ram.memory[80][1] ;
 wire \u_cpu.rf_ram.memory[80][2] ;
 wire \u_cpu.rf_ram.memory[80][3] ;
 wire \u_cpu.rf_ram.memory[80][4] ;
 wire \u_cpu.rf_ram.memory[80][5] ;
 wire \u_cpu.rf_ram.memory[80][6] ;
 wire \u_cpu.rf_ram.memory[80][7] ;
 wire \u_cpu.rf_ram.memory[81][0] ;
 wire \u_cpu.rf_ram.memory[81][1] ;
 wire \u_cpu.rf_ram.memory[81][2] ;
 wire \u_cpu.rf_ram.memory[81][3] ;
 wire \u_cpu.rf_ram.memory[81][4] ;
 wire \u_cpu.rf_ram.memory[81][5] ;
 wire \u_cpu.rf_ram.memory[81][6] ;
 wire \u_cpu.rf_ram.memory[81][7] ;
 wire \u_cpu.rf_ram.memory[82][0] ;
 wire \u_cpu.rf_ram.memory[82][1] ;
 wire \u_cpu.rf_ram.memory[82][2] ;
 wire \u_cpu.rf_ram.memory[82][3] ;
 wire \u_cpu.rf_ram.memory[82][4] ;
 wire \u_cpu.rf_ram.memory[82][5] ;
 wire \u_cpu.rf_ram.memory[82][6] ;
 wire \u_cpu.rf_ram.memory[82][7] ;
 wire \u_cpu.rf_ram.memory[83][0] ;
 wire \u_cpu.rf_ram.memory[83][1] ;
 wire \u_cpu.rf_ram.memory[83][2] ;
 wire \u_cpu.rf_ram.memory[83][3] ;
 wire \u_cpu.rf_ram.memory[83][4] ;
 wire \u_cpu.rf_ram.memory[83][5] ;
 wire \u_cpu.rf_ram.memory[83][6] ;
 wire \u_cpu.rf_ram.memory[83][7] ;
 wire \u_cpu.rf_ram.memory[84][0] ;
 wire \u_cpu.rf_ram.memory[84][1] ;
 wire \u_cpu.rf_ram.memory[84][2] ;
 wire \u_cpu.rf_ram.memory[84][3] ;
 wire \u_cpu.rf_ram.memory[84][4] ;
 wire \u_cpu.rf_ram.memory[84][5] ;
 wire \u_cpu.rf_ram.memory[84][6] ;
 wire \u_cpu.rf_ram.memory[84][7] ;
 wire \u_cpu.rf_ram.memory[85][0] ;
 wire \u_cpu.rf_ram.memory[85][1] ;
 wire \u_cpu.rf_ram.memory[85][2] ;
 wire \u_cpu.rf_ram.memory[85][3] ;
 wire \u_cpu.rf_ram.memory[85][4] ;
 wire \u_cpu.rf_ram.memory[85][5] ;
 wire \u_cpu.rf_ram.memory[85][6] ;
 wire \u_cpu.rf_ram.memory[85][7] ;
 wire \u_cpu.rf_ram.memory[86][0] ;
 wire \u_cpu.rf_ram.memory[86][1] ;
 wire \u_cpu.rf_ram.memory[86][2] ;
 wire \u_cpu.rf_ram.memory[86][3] ;
 wire \u_cpu.rf_ram.memory[86][4] ;
 wire \u_cpu.rf_ram.memory[86][5] ;
 wire \u_cpu.rf_ram.memory[86][6] ;
 wire \u_cpu.rf_ram.memory[86][7] ;
 wire \u_cpu.rf_ram.memory[87][0] ;
 wire \u_cpu.rf_ram.memory[87][1] ;
 wire \u_cpu.rf_ram.memory[87][2] ;
 wire \u_cpu.rf_ram.memory[87][3] ;
 wire \u_cpu.rf_ram.memory[87][4] ;
 wire \u_cpu.rf_ram.memory[87][5] ;
 wire \u_cpu.rf_ram.memory[87][6] ;
 wire \u_cpu.rf_ram.memory[87][7] ;
 wire \u_cpu.rf_ram.memory[88][0] ;
 wire \u_cpu.rf_ram.memory[88][1] ;
 wire \u_cpu.rf_ram.memory[88][2] ;
 wire \u_cpu.rf_ram.memory[88][3] ;
 wire \u_cpu.rf_ram.memory[88][4] ;
 wire \u_cpu.rf_ram.memory[88][5] ;
 wire \u_cpu.rf_ram.memory[88][6] ;
 wire \u_cpu.rf_ram.memory[88][7] ;
 wire \u_cpu.rf_ram.memory[89][0] ;
 wire \u_cpu.rf_ram.memory[89][1] ;
 wire \u_cpu.rf_ram.memory[89][2] ;
 wire \u_cpu.rf_ram.memory[89][3] ;
 wire \u_cpu.rf_ram.memory[89][4] ;
 wire \u_cpu.rf_ram.memory[89][5] ;
 wire \u_cpu.rf_ram.memory[89][6] ;
 wire \u_cpu.rf_ram.memory[89][7] ;
 wire \u_cpu.rf_ram.memory[8][0] ;
 wire \u_cpu.rf_ram.memory[8][1] ;
 wire \u_cpu.rf_ram.memory[8][2] ;
 wire \u_cpu.rf_ram.memory[8][3] ;
 wire \u_cpu.rf_ram.memory[8][4] ;
 wire \u_cpu.rf_ram.memory[8][5] ;
 wire \u_cpu.rf_ram.memory[8][6] ;
 wire \u_cpu.rf_ram.memory[8][7] ;
 wire \u_cpu.rf_ram.memory[90][0] ;
 wire \u_cpu.rf_ram.memory[90][1] ;
 wire \u_cpu.rf_ram.memory[90][2] ;
 wire \u_cpu.rf_ram.memory[90][3] ;
 wire \u_cpu.rf_ram.memory[90][4] ;
 wire \u_cpu.rf_ram.memory[90][5] ;
 wire \u_cpu.rf_ram.memory[90][6] ;
 wire \u_cpu.rf_ram.memory[90][7] ;
 wire \u_cpu.rf_ram.memory[91][0] ;
 wire \u_cpu.rf_ram.memory[91][1] ;
 wire \u_cpu.rf_ram.memory[91][2] ;
 wire \u_cpu.rf_ram.memory[91][3] ;
 wire \u_cpu.rf_ram.memory[91][4] ;
 wire \u_cpu.rf_ram.memory[91][5] ;
 wire \u_cpu.rf_ram.memory[91][6] ;
 wire \u_cpu.rf_ram.memory[91][7] ;
 wire \u_cpu.rf_ram.memory[92][0] ;
 wire \u_cpu.rf_ram.memory[92][1] ;
 wire \u_cpu.rf_ram.memory[92][2] ;
 wire \u_cpu.rf_ram.memory[92][3] ;
 wire \u_cpu.rf_ram.memory[92][4] ;
 wire \u_cpu.rf_ram.memory[92][5] ;
 wire \u_cpu.rf_ram.memory[92][6] ;
 wire \u_cpu.rf_ram.memory[92][7] ;
 wire \u_cpu.rf_ram.memory[93][0] ;
 wire \u_cpu.rf_ram.memory[93][1] ;
 wire \u_cpu.rf_ram.memory[93][2] ;
 wire \u_cpu.rf_ram.memory[93][3] ;
 wire \u_cpu.rf_ram.memory[93][4] ;
 wire \u_cpu.rf_ram.memory[93][5] ;
 wire \u_cpu.rf_ram.memory[93][6] ;
 wire \u_cpu.rf_ram.memory[93][7] ;
 wire \u_cpu.rf_ram.memory[94][0] ;
 wire \u_cpu.rf_ram.memory[94][1] ;
 wire \u_cpu.rf_ram.memory[94][2] ;
 wire \u_cpu.rf_ram.memory[94][3] ;
 wire \u_cpu.rf_ram.memory[94][4] ;
 wire \u_cpu.rf_ram.memory[94][5] ;
 wire \u_cpu.rf_ram.memory[94][6] ;
 wire \u_cpu.rf_ram.memory[94][7] ;
 wire \u_cpu.rf_ram.memory[95][0] ;
 wire \u_cpu.rf_ram.memory[95][1] ;
 wire \u_cpu.rf_ram.memory[95][2] ;
 wire \u_cpu.rf_ram.memory[95][3] ;
 wire \u_cpu.rf_ram.memory[95][4] ;
 wire \u_cpu.rf_ram.memory[95][5] ;
 wire \u_cpu.rf_ram.memory[95][6] ;
 wire \u_cpu.rf_ram.memory[95][7] ;
 wire \u_cpu.rf_ram.memory[96][0] ;
 wire \u_cpu.rf_ram.memory[96][1] ;
 wire \u_cpu.rf_ram.memory[96][2] ;
 wire \u_cpu.rf_ram.memory[96][3] ;
 wire \u_cpu.rf_ram.memory[96][4] ;
 wire \u_cpu.rf_ram.memory[96][5] ;
 wire \u_cpu.rf_ram.memory[96][6] ;
 wire \u_cpu.rf_ram.memory[96][7] ;
 wire \u_cpu.rf_ram.memory[97][0] ;
 wire \u_cpu.rf_ram.memory[97][1] ;
 wire \u_cpu.rf_ram.memory[97][2] ;
 wire \u_cpu.rf_ram.memory[97][3] ;
 wire \u_cpu.rf_ram.memory[97][4] ;
 wire \u_cpu.rf_ram.memory[97][5] ;
 wire \u_cpu.rf_ram.memory[97][6] ;
 wire \u_cpu.rf_ram.memory[97][7] ;
 wire \u_cpu.rf_ram.memory[98][0] ;
 wire \u_cpu.rf_ram.memory[98][1] ;
 wire \u_cpu.rf_ram.memory[98][2] ;
 wire \u_cpu.rf_ram.memory[98][3] ;
 wire \u_cpu.rf_ram.memory[98][4] ;
 wire \u_cpu.rf_ram.memory[98][5] ;
 wire \u_cpu.rf_ram.memory[98][6] ;
 wire \u_cpu.rf_ram.memory[98][7] ;
 wire \u_cpu.rf_ram.memory[99][0] ;
 wire \u_cpu.rf_ram.memory[99][1] ;
 wire \u_cpu.rf_ram.memory[99][2] ;
 wire \u_cpu.rf_ram.memory[99][3] ;
 wire \u_cpu.rf_ram.memory[99][4] ;
 wire \u_cpu.rf_ram.memory[99][5] ;
 wire \u_cpu.rf_ram.memory[99][6] ;
 wire \u_cpu.rf_ram.memory[99][7] ;
 wire \u_cpu.rf_ram.memory[9][0] ;
 wire \u_cpu.rf_ram.memory[9][1] ;
 wire \u_cpu.rf_ram.memory[9][2] ;
 wire \u_cpu.rf_ram.memory[9][3] ;
 wire \u_cpu.rf_ram.memory[9][4] ;
 wire \u_cpu.rf_ram.memory[9][5] ;
 wire \u_cpu.rf_ram.memory[9][6] ;
 wire \u_cpu.rf_ram.memory[9][7] ;
 wire \u_cpu.rf_ram.rdata[0] ;
 wire \u_cpu.rf_ram.rdata[1] ;
 wire \u_cpu.rf_ram.rdata[2] ;
 wire \u_cpu.rf_ram.rdata[3] ;
 wire \u_cpu.rf_ram.rdata[4] ;
 wire \u_cpu.rf_ram.rdata[5] ;
 wire \u_cpu.rf_ram.rdata[6] ;
 wire \u_cpu.rf_ram.rdata[7] ;
 wire \u_cpu.rf_ram.regzero ;
 wire \u_cpu.rf_ram_if.genblk1.wtrig0_r ;
 wire \u_cpu.rf_ram_if.rcnt[0] ;
 wire \u_cpu.rf_ram_if.rcnt[1] ;
 wire \u_cpu.rf_ram_if.rcnt[2] ;
 wire \u_cpu.rf_ram_if.rdata0[1] ;
 wire \u_cpu.rf_ram_if.rdata0[2] ;
 wire \u_cpu.rf_ram_if.rdata0[3] ;
 wire \u_cpu.rf_ram_if.rdata0[4] ;
 wire \u_cpu.rf_ram_if.rdata0[5] ;
 wire \u_cpu.rf_ram_if.rdata0[6] ;
 wire \u_cpu.rf_ram_if.rdata0[7] ;
 wire \u_cpu.rf_ram_if.rdata1[0] ;
 wire \u_cpu.rf_ram_if.rdata1[1] ;
 wire \u_cpu.rf_ram_if.rdata1[2] ;
 wire \u_cpu.rf_ram_if.rdata1[3] ;
 wire \u_cpu.rf_ram_if.rdata1[4] ;
 wire \u_cpu.rf_ram_if.rdata1[5] ;
 wire \u_cpu.rf_ram_if.rdata1[6] ;
 wire \u_cpu.rf_ram_if.rgnt ;
 wire \u_cpu.rf_ram_if.rreq_r ;
 wire \u_cpu.rf_ram_if.rtrig0 ;
 wire \u_cpu.rf_ram_if.rtrig1 ;
 wire \u_cpu.rf_ram_if.wdata0_r[0] ;
 wire \u_cpu.rf_ram_if.wdata0_r[1] ;
 wire \u_cpu.rf_ram_if.wdata0_r[2] ;
 wire \u_cpu.rf_ram_if.wdata0_r[3] ;
 wire \u_cpu.rf_ram_if.wdata0_r[4] ;
 wire \u_cpu.rf_ram_if.wdata0_r[5] ;
 wire \u_cpu.rf_ram_if.wdata0_r[6] ;
 wire \u_cpu.rf_ram_if.wdata1_r[0] ;
 wire \u_cpu.rf_ram_if.wdata1_r[1] ;
 wire \u_cpu.rf_ram_if.wdata1_r[2] ;
 wire \u_cpu.rf_ram_if.wdata1_r[3] ;
 wire \u_cpu.rf_ram_if.wdata1_r[4] ;
 wire \u_cpu.rf_ram_if.wdata1_r[5] ;
 wire \u_cpu.rf_ram_if.wdata1_r[6] ;
 wire \u_cpu.rf_ram_if.wdata1_r[7] ;
 wire \u_cpu.rf_ram_if.wen0_r ;
 wire \u_cpu.rf_ram_if.wen1_r ;
 wire \u_cpu.rf_ram_if.wtrig0 ;
 wire \u_scanchain_local.clk ;
 wire \u_scanchain_local.clk_out ;
 wire \u_scanchain_local.data_out ;
 wire \u_scanchain_local.data_out_i ;
 wire \u_scanchain_local.module_data_in[34] ;
 wire \u_scanchain_local.module_data_in[35] ;
 wire \u_scanchain_local.module_data_in[36] ;
 wire \u_scanchain_local.module_data_in[37] ;
 wire \u_scanchain_local.module_data_in[38] ;
 wire \u_scanchain_local.module_data_in[39] ;
 wire \u_scanchain_local.module_data_in[40] ;
 wire \u_scanchain_local.module_data_in[41] ;
 wire \u_scanchain_local.module_data_in[42] ;
 wire \u_scanchain_local.module_data_in[43] ;
 wire \u_scanchain_local.module_data_in[44] ;
 wire \u_scanchain_local.module_data_in[45] ;
 wire \u_scanchain_local.module_data_in[46] ;
 wire \u_scanchain_local.module_data_in[47] ;
 wire \u_scanchain_local.module_data_in[48] ;
 wire \u_scanchain_local.module_data_in[49] ;
 wire \u_scanchain_local.module_data_in[50] ;
 wire \u_scanchain_local.module_data_in[51] ;
 wire \u_scanchain_local.module_data_in[52] ;
 wire \u_scanchain_local.module_data_in[53] ;
 wire \u_scanchain_local.module_data_in[54] ;
 wire \u_scanchain_local.module_data_in[55] ;
 wire \u_scanchain_local.module_data_in[56] ;
 wire \u_scanchain_local.module_data_in[57] ;
 wire \u_scanchain_local.module_data_in[58] ;
 wire \u_scanchain_local.module_data_in[59] ;
 wire \u_scanchain_local.module_data_in[60] ;
 wire \u_scanchain_local.module_data_in[61] ;
 wire \u_scanchain_local.module_data_in[62] ;
 wire \u_scanchain_local.module_data_in[63] ;
 wire \u_scanchain_local.module_data_in[64] ;
 wire \u_scanchain_local.module_data_in[65] ;
 wire \u_scanchain_local.module_data_in[66] ;
 wire \u_scanchain_local.module_data_in[67] ;
 wire \u_scanchain_local.module_data_in[68] ;
 wire \u_scanchain_local.module_data_in[69] ;

 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _04838_ (.I(\u_cpu.rf_ram_if.rcnt[0] ),
    .ZN(_01366_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _04839_ (.A1(\u_cpu.rf_ram_if.rcnt[2] ),
    .A2(\u_cpu.rf_ram_if.rcnt[1] ),
    .A3(_01366_),
    .Z(_01367_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _04840_ (.I(_01367_),
    .Z(_01368_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _04841_ (.I(_01368_),
    .ZN(\u_cpu.rf_ram_if.rtrig0 ));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _04842_ (.A1(\u_cpu.cpu.bufreg.lsb[0] ),
    .A2(\u_cpu.cpu.bufreg.lsb[1] ),
    .ZN(\u_arbiter.i_wb_cpu_dbus_sel[0] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _04843_ (.I(\u_cpu.cpu.csr_d_sel ),
    .Z(_01369_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _04844_ (.I(\u_cpu.cpu.decode.co_mem_word ),
    .Z(_01370_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _04845_ (.A1(_01369_),
    .A2(_01370_),
    .A3(\u_cpu.cpu.bne_or_bge ),
    .ZN(_01371_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _04846_ (.I(\u_cpu.cpu.decode.opcode[2] ),
    .Z(_01372_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _04847_ (.I(_01372_),
    .ZN(_01373_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _04848_ (.I(\u_cpu.cpu.branch_op ),
    .Z(_01374_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _04849_ (.I(_01374_),
    .ZN(_01375_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _04850_ (.A1(_01373_),
    .A2(_01375_),
    .ZN(_01376_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _04851_ (.A1(\u_cpu.cpu.decode.op21 ),
    .A2(_01371_),
    .A3(_01376_),
    .ZN(_01377_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _04852_ (.A1(_01372_),
    .A2(_01374_),
    .ZN(_01378_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _04853_ (.A1(_01371_),
    .A2(_01378_),
    .ZN(_01379_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _04854_ (.I(\u_cpu.cpu.decode.op26 ),
    .ZN(_01380_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _04855_ (.I(\u_cpu.cpu.decode.co_ebreak ),
    .ZN(_01381_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _04856_ (.A1(\u_cpu.cpu.decode.op21 ),
    .A2(_01380_),
    .B(_01381_),
    .ZN(_01382_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _04857_ (.A1(_01369_),
    .A2(_01370_),
    .A3(\u_cpu.cpu.decode.op21 ),
    .A4(\u_cpu.cpu.bne_or_bge ),
    .Z(_01383_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _04858_ (.I(\u_cpu.cpu.genblk3.csr.o_new_irq ),
    .ZN(_01384_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _04859_ (.I(\u_cpu.cpu.state.genblk1.misalign_trap_sync_r ),
    .ZN(_01385_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _04860_ (.A1(_01378_),
    .A2(_01383_),
    .B(_01384_),
    .C(_01385_),
    .ZN(_01386_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _04861_ (.A1(_01379_),
    .A2(_01382_),
    .B(_01386_),
    .ZN(_01387_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _04862_ (.A1(\u_cpu.rf_ram_if.rtrig0 ),
    .A2(_01377_),
    .A3(_01387_),
    .Z(_01388_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _04863_ (.A1(\u_cpu.cpu.immdec.imm24_20[0] ),
    .A2(_01388_),
    .Z(_01389_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _04864_ (.I(\u_cpu.cpu.csr_imm ),
    .ZN(_01390_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _04865_ (.A1(_01390_),
    .A2(\u_cpu.rf_ram_if.rtrig0 ),
    .ZN(_01391_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _04866_ (.A1(_01378_),
    .A2(_01383_),
    .ZN(_01392_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _04867_ (.A1(\u_cpu.cpu.genblk3.csr.o_new_irq ),
    .A2(\u_cpu.cpu.state.genblk1.misalign_trap_sync_r ),
    .A3(_01392_),
    .ZN(_01393_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _04868_ (.A1(\u_cpu.cpu.decode.op21 ),
    .A2(_01380_),
    .ZN(_01394_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _04869_ (.A1(_01393_),
    .A2(_01394_),
    .B(_01387_),
    .C(_01368_),
    .ZN(_01395_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _04870_ (.A1(_01389_),
    .A2(_01391_),
    .A3(_01395_),
    .Z(_01396_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _04871_ (.I(_01396_),
    .Z(_01397_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _04872_ (.I(_01397_),
    .Z(_01398_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _04873_ (.I(_01398_),
    .Z(_01399_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _04874_ (.A1(\u_cpu.cpu.immdec.imm19_12_20[8] ),
    .A2(_01368_),
    .ZN(_01400_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _04875_ (.A1(\u_cpu.cpu.immdec.imm24_20[4] ),
    .A2(_01388_),
    .ZN(_01401_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _04876_ (.A1(_01400_),
    .A2(_01401_),
    .ZN(_01402_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _04877_ (.I(_01368_),
    .Z(_01403_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _04878_ (.A1(_01377_),
    .A2(_01387_),
    .B(_01403_),
    .ZN(_01404_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _04879_ (.A1(_01402_),
    .A2(_01404_),
    .ZN(_01405_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _04880_ (.I(_01405_),
    .Z(_01406_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _04881_ (.A1(\u_cpu.cpu.immdec.imm19_12_20[5] ),
    .A2(\u_cpu.rf_ram_if.rtrig0 ),
    .ZN(_01407_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _04882_ (.I(_01369_),
    .ZN(_01408_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _04883_ (.A1(_01370_),
    .A2(\u_cpu.cpu.bne_or_bge ),
    .ZN(_01409_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _04884_ (.A1(_01408_),
    .A2(_01409_),
    .ZN(_01410_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _04885_ (.A1(_01410_),
    .A2(_01376_),
    .ZN(_01411_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _04886_ (.A1(\u_cpu.cpu.decode.op26 ),
    .A2(\u_cpu.cpu.decode.co_ebreak ),
    .ZN(_01412_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _04887_ (.A1(_01411_),
    .A2(_01412_),
    .B(\u_cpu.rf_ram_if.rtrig0 ),
    .C(_01377_),
    .ZN(_01413_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _04888_ (.A1(\u_cpu.cpu.immdec.imm24_20[1] ),
    .A2(_01387_),
    .B(_01413_),
    .ZN(_01414_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _04889_ (.A1(_01407_),
    .A2(_01414_),
    .Z(_01415_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _04890_ (.I(_01415_),
    .Z(_01416_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _04891_ (.I(_01416_),
    .Z(_01417_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _04892_ (.I(_01417_),
    .Z(_01418_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _04893_ (.A1(\u_cpu.cpu.immdec.imm19_12_20[7] ),
    .A2(_01368_),
    .ZN(_01419_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _04894_ (.A1(\u_cpu.cpu.immdec.imm24_20[3] ),
    .A2(_01388_),
    .ZN(_01420_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _04895_ (.A1(_01419_),
    .A2(_01420_),
    .Z(_01421_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _04896_ (.I(_01421_),
    .Z(_01422_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _04897_ (.A1(\u_cpu.cpu.immdec.imm19_12_20[6] ),
    .A2(_01368_),
    .ZN(_01423_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _04898_ (.A1(\u_cpu.cpu.immdec.imm24_20[2] ),
    .A2(_01388_),
    .ZN(_01424_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _04899_ (.A1(_01423_),
    .A2(_01424_),
    .Z(_01425_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _04900_ (.I(_01425_),
    .Z(_01426_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _04901_ (.A1(_01406_),
    .A2(_01418_),
    .A3(_01422_),
    .A4(_01426_),
    .ZN(_01427_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _04902_ (.A1(_01399_),
    .A2(_01427_),
    .ZN(_00025_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _04903_ (.I(_01403_),
    .ZN(\u_cpu.rf_ram_if.wtrig0 ));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _04904_ (.I(io_in[1]),
    .Z(_01428_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _04905_ (.I(_01428_),
    .ZN(_01429_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _04906_ (.A1(_01429_),
    .A2(\u_cpu.cpu.state.ibus_cyc ),
    .Z(_01430_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _04907_ (.I(_01430_),
    .Z(_01431_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _04908_ (.A1(\u_arbiter.i_wb_cpu_ibus_adr[0] ),
    .A2(_01431_),
    .Z(_01432_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _04909_ (.I(_01432_),
    .Z(\u_arbiter.o_wb_cpu_adr[0] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _04910_ (.A1(\u_arbiter.i_wb_cpu_ibus_adr[1] ),
    .A2(_01431_),
    .Z(_01433_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _04911_ (.I(_01433_),
    .Z(\u_arbiter.o_wb_cpu_adr[1] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _04912_ (.I(\u_cpu.cpu.genblk1.align.ctrl_misal ),
    .Z(_01434_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _04913_ (.I(_01434_),
    .Z(_01435_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _04914_ (.I(_01435_),
    .Z(_01436_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _04915_ (.I(_01436_),
    .Z(_01437_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _04916_ (.A1(_01437_),
    .A2(\u_cpu.cpu.ctrl.o_ibus_adr[2] ),
    .ZN(_01438_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _04917_ (.A1(_01437_),
    .A2(\u_cpu.cpu.ctrl.o_ibus_adr[2] ),
    .ZN(_01439_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _04918_ (.A1(_01431_),
    .A2(_01439_),
    .ZN(_01440_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _04919_ (.A1(_01429_),
    .A2(\u_cpu.cpu.state.ibus_cyc ),
    .ZN(_01441_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _04920_ (.I(_01441_),
    .Z(_01442_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _04921_ (.I(_01442_),
    .Z(_01443_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _04922_ (.A1(\u_arbiter.i_wb_cpu_dbus_adr[2] ),
    .A2(_01443_),
    .ZN(_01444_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _04923_ (.A1(_01438_),
    .A2(_01440_),
    .B(_01444_),
    .ZN(\u_arbiter.o_wb_cpu_adr[2] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _04924_ (.I(_01442_),
    .Z(_01445_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _04925_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[3] ),
    .A2(_01439_),
    .Z(_01446_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _04926_ (.A1(\u_arbiter.i_wb_cpu_dbus_adr[3] ),
    .A2(_01443_),
    .ZN(_01447_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _04927_ (.A1(_01445_),
    .A2(_01446_),
    .B(_01447_),
    .ZN(\u_arbiter.o_wb_cpu_adr[3] ));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _04928_ (.A1(_01437_),
    .A2(\u_cpu.cpu.ctrl.o_ibus_adr[3] ),
    .A3(\u_cpu.cpu.ctrl.o_ibus_adr[2] ),
    .ZN(_01448_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _04929_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[4] ),
    .A2(_01448_),
    .Z(_01449_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _04930_ (.A1(\u_arbiter.i_wb_cpu_dbus_adr[4] ),
    .A2(_01443_),
    .ZN(_01450_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _04931_ (.A1(_01445_),
    .A2(_01449_),
    .B(_01450_),
    .ZN(\u_arbiter.o_wb_cpu_adr[4] ));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _04932_ (.A1(_01434_),
    .A2(\u_cpu.cpu.ctrl.o_ibus_adr[4] ),
    .A3(\u_cpu.cpu.ctrl.o_ibus_adr[3] ),
    .A4(\u_cpu.cpu.ctrl.o_ibus_adr[2] ),
    .Z(_01451_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _04933_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[5] ),
    .A2(_01451_),
    .ZN(_01452_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _04934_ (.A1(\u_arbiter.i_wb_cpu_dbus_adr[5] ),
    .A2(_01443_),
    .ZN(_01453_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _04935_ (.A1(_01445_),
    .A2(_01452_),
    .B(_01453_),
    .ZN(\u_arbiter.o_wb_cpu_adr[5] ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _04936_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[5] ),
    .A2(_01451_),
    .B(\u_cpu.cpu.ctrl.o_ibus_adr[6] ),
    .ZN(_01454_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _04937_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[6] ),
    .A2(\u_cpu.cpu.ctrl.o_ibus_adr[5] ),
    .A3(_01451_),
    .ZN(_01455_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _04938_ (.A1(_01431_),
    .A2(_01455_),
    .ZN(_01456_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _04939_ (.I(_01442_),
    .Z(_01457_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _04940_ (.A1(\u_arbiter.i_wb_cpu_dbus_adr[6] ),
    .A2(_01457_),
    .ZN(_01458_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _04941_ (.A1(_01454_),
    .A2(_01456_),
    .B(_01458_),
    .ZN(\u_arbiter.o_wb_cpu_adr[6] ));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _04942_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[7] ),
    .A2(_01455_),
    .Z(_01459_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _04943_ (.A1(\u_arbiter.i_wb_cpu_dbus_adr[7] ),
    .A2(_01457_),
    .ZN(_01460_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _04944_ (.A1(_01445_),
    .A2(_01459_),
    .B(_01460_),
    .ZN(\u_arbiter.o_wb_cpu_adr[7] ));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _04945_ (.I(\u_cpu.cpu.ctrl.o_ibus_adr[8] ),
    .ZN(_01461_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _04946_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[7] ),
    .A2(\u_cpu.cpu.ctrl.o_ibus_adr[6] ),
    .A3(\u_cpu.cpu.ctrl.o_ibus_adr[5] ),
    .A4(_01451_),
    .ZN(_01462_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _04947_ (.A1(_01461_),
    .A2(_01462_),
    .ZN(_01463_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _04948_ (.A1(_01461_),
    .A2(_01462_),
    .Z(_01464_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _04949_ (.A1(_01463_),
    .A2(_01464_),
    .ZN(_01465_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _04950_ (.A1(\u_arbiter.i_wb_cpu_dbus_adr[8] ),
    .A2(_01457_),
    .ZN(_01466_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _04951_ (.A1(_01445_),
    .A2(_01465_),
    .B(_01466_),
    .ZN(\u_arbiter.o_wb_cpu_adr[8] ));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _04952_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[9] ),
    .A2(_01464_),
    .Z(_01467_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _04953_ (.A1(\u_arbiter.i_wb_cpu_dbus_adr[9] ),
    .A2(_01457_),
    .ZN(_01468_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _04954_ (.A1(_01445_),
    .A2(_01467_),
    .B(_01468_),
    .ZN(\u_arbiter.o_wb_cpu_adr[9] ));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _04955_ (.A1(\u_arbiter.i_wb_cpu_dbus_adr[10] ),
    .A2(_01443_),
    .ZN(_01469_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _04956_ (.I(\u_cpu.cpu.ctrl.o_ibus_adr[9] ),
    .ZN(_01470_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _04957_ (.A1(_01470_),
    .A2(_01464_),
    .ZN(_01471_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _04958_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[10] ),
    .A2(_01471_),
    .B(_01442_),
    .ZN(_01472_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _04959_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[10] ),
    .A2(_01471_),
    .B(_01472_),
    .ZN(_01473_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _04960_ (.A1(_01469_),
    .A2(_01473_),
    .ZN(\u_arbiter.o_wb_cpu_adr[10] ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _04961_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[10] ),
    .A2(_01471_),
    .B(\u_cpu.cpu.ctrl.o_ibus_adr[11] ),
    .ZN(_01474_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _04962_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[11] ),
    .A2(\u_cpu.cpu.ctrl.o_ibus_adr[10] ),
    .ZN(_01475_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _04963_ (.A1(_01470_),
    .A2(_01461_),
    .A3(_01462_),
    .A4(_01475_),
    .ZN(_01476_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _04964_ (.A1(\u_arbiter.i_wb_cpu_dbus_adr[11] ),
    .A2(_01457_),
    .ZN(_01477_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _04965_ (.A1(_01443_),
    .A2(_01474_),
    .A3(_01476_),
    .B(_01477_),
    .ZN(\u_arbiter.o_wb_cpu_adr[11] ));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _04966_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[12] ),
    .A2(_01476_),
    .ZN(_01478_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _04967_ (.A1(\u_arbiter.i_wb_cpu_dbus_adr[12] ),
    .A2(_01457_),
    .ZN(_01479_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _04968_ (.A1(_01445_),
    .A2(_01478_),
    .B(_01479_),
    .ZN(\u_arbiter.o_wb_cpu_adr[12] ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _04969_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[12] ),
    .A2(_01476_),
    .B(\u_cpu.cpu.ctrl.o_ibus_adr[13] ),
    .ZN(_01480_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _04970_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[13] ),
    .A2(\u_cpu.cpu.ctrl.o_ibus_adr[12] ),
    .A3(_01476_),
    .Z(_01481_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _04971_ (.A1(\u_arbiter.i_wb_cpu_dbus_adr[13] ),
    .A2(_01442_),
    .ZN(_01482_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _04972_ (.A1(_01443_),
    .A2(_01480_),
    .A3(_01481_),
    .B(_01482_),
    .ZN(\u_arbiter.o_wb_cpu_adr[13] ));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _04973_ (.A1(\u_arbiter.i_wb_cpu_dbus_adr[14] ),
    .A2(_01443_),
    .ZN(_01483_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _04974_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[14] ),
    .A2(_01481_),
    .B(_01442_),
    .ZN(_01484_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _04975_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[14] ),
    .A2(_01481_),
    .B(_01484_),
    .ZN(_01485_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _04976_ (.A1(_01483_),
    .A2(_01485_),
    .ZN(\u_arbiter.o_wb_cpu_adr[14] ));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _04977_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[14] ),
    .A2(_01481_),
    .B(\u_cpu.cpu.ctrl.o_ibus_adr[15] ),
    .ZN(_01486_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _04978_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[15] ),
    .A2(\u_cpu.cpu.ctrl.o_ibus_adr[14] ),
    .Z(_01487_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _04979_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[13] ),
    .A2(\u_cpu.cpu.ctrl.o_ibus_adr[12] ),
    .A3(_01476_),
    .A4(_01487_),
    .Z(_01488_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _04980_ (.A1(\u_arbiter.i_wb_cpu_dbus_adr[15] ),
    .A2(_01442_),
    .ZN(_01489_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _04981_ (.A1(_01443_),
    .A2(_01486_),
    .A3(_01488_),
    .B(_01489_),
    .ZN(\u_arbiter.o_wb_cpu_adr[15] ));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _04982_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[16] ),
    .A2(_01488_),
    .ZN(_01490_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _04983_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[16] ),
    .A2(_01488_),
    .Z(_01491_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _04984_ (.A1(\u_arbiter.i_wb_cpu_dbus_adr[16] ),
    .A2(_01442_),
    .ZN(_01492_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _04985_ (.A1(_01443_),
    .A2(_01490_),
    .A3(_01491_),
    .B(_01492_),
    .ZN(\u_arbiter.o_wb_cpu_adr[16] ));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _04986_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[17] ),
    .A2(_01491_),
    .ZN(_01493_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _04987_ (.A1(\u_arbiter.i_wb_cpu_dbus_adr[17] ),
    .A2(_01457_),
    .ZN(_01494_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _04988_ (.A1(_01445_),
    .A2(_01493_),
    .B(_01494_),
    .ZN(\u_arbiter.o_wb_cpu_adr[17] ));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _04989_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[18] ),
    .A2(\u_cpu.cpu.ctrl.o_ibus_adr[17] ),
    .A3(\u_cpu.cpu.ctrl.o_ibus_adr[16] ),
    .A4(_01488_),
    .Z(_01495_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _04990_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[17] ),
    .A2(_01491_),
    .B(\u_cpu.cpu.ctrl.o_ibus_adr[18] ),
    .ZN(_01496_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _04991_ (.A1(\u_arbiter.i_wb_cpu_dbus_adr[18] ),
    .A2(_01442_),
    .ZN(_01497_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _04992_ (.A1(_01443_),
    .A2(_01495_),
    .A3(_01496_),
    .B(_01497_),
    .ZN(\u_arbiter.o_wb_cpu_adr[18] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _04993_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[19] ),
    .A2(_01495_),
    .Z(_01498_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _04994_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[19] ),
    .A2(_01495_),
    .ZN(_01499_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _04995_ (.A1(\u_arbiter.i_wb_cpu_dbus_adr[19] ),
    .A2(_01442_),
    .ZN(_01500_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _04996_ (.A1(_01443_),
    .A2(_01498_),
    .A3(_01499_),
    .B(_01500_),
    .ZN(\u_arbiter.o_wb_cpu_adr[19] ));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _04997_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[20] ),
    .A2(_01498_),
    .ZN(_01501_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _04998_ (.A1(\u_arbiter.i_wb_cpu_dbus_adr[20] ),
    .A2(_01457_),
    .ZN(_01502_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _04999_ (.A1(_01445_),
    .A2(_01501_),
    .B(_01502_),
    .ZN(\u_arbiter.o_wb_cpu_adr[20] ));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05000_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[20] ),
    .A2(_01498_),
    .ZN(_01503_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _05001_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[21] ),
    .A2(_01503_),
    .Z(_01504_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05002_ (.A1(\u_arbiter.i_wb_cpu_dbus_adr[21] ),
    .A2(_01457_),
    .ZN(_01505_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05003_ (.A1(_01445_),
    .A2(_01504_),
    .B(_01505_),
    .ZN(\u_arbiter.o_wb_cpu_adr[21] ));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05004_ (.I(\u_cpu.cpu.ctrl.o_ibus_adr[22] ),
    .ZN(_01506_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _05005_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[21] ),
    .A2(\u_cpu.cpu.ctrl.o_ibus_adr[20] ),
    .A3(\u_cpu.cpu.ctrl.o_ibus_adr[19] ),
    .A4(_01495_),
    .ZN(_01507_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _05006_ (.A1(_01506_),
    .A2(_01507_),
    .Z(_01508_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05007_ (.A1(_01506_),
    .A2(_01507_),
    .ZN(_01509_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05008_ (.A1(\u_arbiter.i_wb_cpu_dbus_adr[22] ),
    .A2(_01442_),
    .ZN(_01510_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _05009_ (.A1(_01443_),
    .A2(_01508_),
    .A3(_01509_),
    .B(_01510_),
    .ZN(\u_arbiter.o_wb_cpu_adr[22] ));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05010_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[23] ),
    .A2(_01509_),
    .ZN(_01511_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05011_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[23] ),
    .A2(\u_cpu.cpu.ctrl.o_ibus_adr[22] ),
    .ZN(_01512_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05012_ (.A1(_01507_),
    .A2(_01512_),
    .ZN(_01513_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05013_ (.A1(\u_arbiter.i_wb_cpu_dbus_adr[23] ),
    .A2(_01442_),
    .ZN(_01514_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _05014_ (.A1(_01443_),
    .A2(_01511_),
    .A3(_01513_),
    .B(_01514_),
    .ZN(\u_arbiter.o_wb_cpu_adr[23] ));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _05015_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[24] ),
    .A2(_01513_),
    .ZN(_01515_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05016_ (.A1(\u_arbiter.i_wb_cpu_dbus_adr[24] ),
    .A2(_01457_),
    .ZN(_01516_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05017_ (.A1(_01445_),
    .A2(_01515_),
    .B(_01516_),
    .ZN(\u_arbiter.o_wb_cpu_adr[24] ));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05018_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[24] ),
    .A2(_01513_),
    .ZN(_01517_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _05019_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[25] ),
    .A2(_01517_),
    .Z(_01518_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05020_ (.A1(\u_arbiter.i_wb_cpu_dbus_adr[25] ),
    .A2(_01457_),
    .ZN(_01519_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05021_ (.A1(_01445_),
    .A2(_01518_),
    .B(_01519_),
    .ZN(\u_arbiter.o_wb_cpu_adr[25] ));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _05022_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[25] ),
    .A2(\u_cpu.cpu.ctrl.o_ibus_adr[24] ),
    .A3(_01513_),
    .ZN(_01520_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _05023_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[26] ),
    .A2(_01520_),
    .Z(_01521_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05024_ (.A1(\u_arbiter.i_wb_cpu_dbus_adr[26] ),
    .A2(_01457_),
    .ZN(_01522_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05025_ (.A1(_01445_),
    .A2(_01521_),
    .B(_01522_),
    .ZN(\u_arbiter.o_wb_cpu_adr[26] ));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _05026_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[26] ),
    .A2(\u_cpu.cpu.ctrl.o_ibus_adr[25] ),
    .A3(\u_cpu.cpu.ctrl.o_ibus_adr[24] ),
    .A4(_01513_),
    .Z(_01523_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _05027_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[27] ),
    .A2(_01523_),
    .ZN(_01524_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05028_ (.A1(\u_arbiter.i_wb_cpu_dbus_adr[27] ),
    .A2(_01457_),
    .ZN(_01525_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05029_ (.A1(_01445_),
    .A2(_01524_),
    .B(_01525_),
    .ZN(\u_arbiter.o_wb_cpu_adr[27] ));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05030_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[27] ),
    .A2(_01523_),
    .ZN(_01526_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _05031_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[28] ),
    .A2(_01526_),
    .Z(_01527_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05032_ (.A1(\u_arbiter.i_wb_cpu_dbus_adr[28] ),
    .A2(_01457_),
    .ZN(_01528_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05033_ (.A1(_01445_),
    .A2(_01527_),
    .B(_01528_),
    .ZN(\u_arbiter.o_wb_cpu_adr[28] ));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _05034_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[28] ),
    .A2(\u_cpu.cpu.ctrl.o_ibus_adr[27] ),
    .A3(_01523_),
    .ZN(_01529_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _05035_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[29] ),
    .A2(_01529_),
    .Z(_01530_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05036_ (.A1(\u_arbiter.i_wb_cpu_dbus_adr[29] ),
    .A2(_01457_),
    .ZN(_01531_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05037_ (.A1(_01443_),
    .A2(_01530_),
    .B(_01531_),
    .ZN(\u_arbiter.o_wb_cpu_adr[29] ));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _05038_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[29] ),
    .A2(\u_cpu.cpu.ctrl.o_ibus_adr[28] ),
    .A3(\u_cpu.cpu.ctrl.o_ibus_adr[27] ),
    .A4(_01523_),
    .ZN(_01532_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _05039_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[30] ),
    .A2(_01532_),
    .Z(_01533_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05040_ (.A1(\u_arbiter.i_wb_cpu_dbus_adr[30] ),
    .A2(_01457_),
    .ZN(_01534_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05041_ (.A1(_01443_),
    .A2(_01533_),
    .B(_01534_),
    .ZN(\u_arbiter.o_wb_cpu_adr[30] ));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05042_ (.I(\u_cpu.cpu.ctrl.o_ibus_adr[30] ),
    .ZN(_01535_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05043_ (.A1(_01535_),
    .A2(_01532_),
    .ZN(_01536_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _05044_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[31] ),
    .A2(_01536_),
    .Z(_01537_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05045_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[31] ),
    .I1(_01537_),
    .S(_01431_),
    .Z(_01538_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05046_ (.I(_01538_),
    .Z(\u_arbiter.o_wb_cpu_adr[31] ));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05047_ (.A1(_01419_),
    .A2(_01420_),
    .ZN(_01539_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _05048_ (.A1(_01389_),
    .A2(_01391_),
    .A3(_01395_),
    .ZN(_01540_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05049_ (.I(_01540_),
    .Z(_01541_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05050_ (.I(_01541_),
    .Z(_01542_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05051_ (.I(\u_cpu.raddr[0] ),
    .Z(_01543_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05052_ (.I(_01543_),
    .Z(_01544_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05053_ (.I(_01544_),
    .Z(_01545_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05054_ (.I(_01545_),
    .Z(_01546_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05055_ (.I(\u_cpu.raddr[1] ),
    .Z(_01547_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05056_ (.I(_01547_),
    .Z(_01548_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05057_ (.I(_01548_),
    .Z(_01549_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05058_ (.I(_01549_),
    .Z(_01550_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05059_ (.I0(\u_cpu.rf_ram.memory[8][0] ),
    .I1(\u_cpu.rf_ram.memory[9][0] ),
    .I2(\u_cpu.rf_ram.memory[10][0] ),
    .I3(\u_cpu.rf_ram.memory[11][0] ),
    .S0(_01546_),
    .S1(_01550_),
    .Z(_01551_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05060_ (.A1(_01542_),
    .A2(_01551_),
    .ZN(_01552_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05061_ (.I(_01397_),
    .Z(_01553_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05062_ (.I(_01553_),
    .Z(_01554_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05063_ (.I(_01543_),
    .Z(_01555_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05064_ (.I(_01555_),
    .Z(_01556_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05065_ (.I(_01548_),
    .Z(_01557_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05066_ (.I0(\u_cpu.rf_ram.memory[12][0] ),
    .I1(\u_cpu.rf_ram.memory[13][0] ),
    .I2(\u_cpu.rf_ram.memory[14][0] ),
    .I3(\u_cpu.rf_ram.memory[15][0] ),
    .S0(_01556_),
    .S1(_01557_),
    .Z(_01558_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05067_ (.A1(_01554_),
    .A2(_01558_),
    .B(_01417_),
    .ZN(_01559_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05068_ (.I0(\u_cpu.rf_ram.memory[4][0] ),
    .I1(\u_cpu.rf_ram.memory[5][0] ),
    .I2(\u_cpu.rf_ram.memory[6][0] ),
    .I3(\u_cpu.rf_ram.memory[7][0] ),
    .S0(_01546_),
    .S1(_01550_),
    .Z(_01560_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05069_ (.A1(_01554_),
    .A2(_01560_),
    .ZN(_01561_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05070_ (.I(_01541_),
    .Z(_01562_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05071_ (.I0(\u_cpu.rf_ram.memory[0][0] ),
    .I1(\u_cpu.rf_ram.memory[1][0] ),
    .I2(\u_cpu.rf_ram.memory[2][0] ),
    .I3(\u_cpu.rf_ram.memory[3][0] ),
    .S0(_01556_),
    .S1(_01557_),
    .Z(_01563_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05072_ (.A1(_01407_),
    .A2(_01414_),
    .ZN(_01564_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05073_ (.I(_01564_),
    .Z(_01565_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05074_ (.A1(_01562_),
    .A2(_01563_),
    .B(_01565_),
    .ZN(_01566_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05075_ (.A1(_01423_),
    .A2(_01424_),
    .ZN(_01567_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05076_ (.I(_01567_),
    .Z(_01568_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _05077_ (.A1(_01552_),
    .A2(_01559_),
    .B1(_01561_),
    .B2(_01566_),
    .C(_01568_),
    .ZN(_01569_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05078_ (.I(_01398_),
    .Z(_01570_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05079_ (.I(_01544_),
    .Z(_01571_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05080_ (.I(_01571_),
    .Z(_01572_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05081_ (.I(_01548_),
    .Z(_01573_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05082_ (.I(_01573_),
    .Z(_01574_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05083_ (.I0(\u_cpu.rf_ram.memory[20][0] ),
    .I1(\u_cpu.rf_ram.memory[21][0] ),
    .I2(\u_cpu.rf_ram.memory[22][0] ),
    .I3(\u_cpu.rf_ram.memory[23][0] ),
    .S0(_01572_),
    .S1(_01574_),
    .Z(_01575_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05084_ (.A1(_01570_),
    .A2(_01575_),
    .ZN(_01576_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05085_ (.I(_01543_),
    .Z(_01577_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05086_ (.I(_01577_),
    .Z(_01578_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05087_ (.I(_01547_),
    .Z(_01579_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05088_ (.I(_01579_),
    .Z(_01580_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05089_ (.I0(\u_cpu.rf_ram.memory[16][0] ),
    .I1(\u_cpu.rf_ram.memory[17][0] ),
    .I2(\u_cpu.rf_ram.memory[18][0] ),
    .I3(\u_cpu.rf_ram.memory[19][0] ),
    .S0(_01578_),
    .S1(_01580_),
    .Z(_01581_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05090_ (.I(_01565_),
    .Z(_01582_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05091_ (.A1(_01562_),
    .A2(_01581_),
    .B(_01582_),
    .ZN(_01583_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05092_ (.I0(\u_cpu.rf_ram.memory[28][0] ),
    .I1(\u_cpu.rf_ram.memory[29][0] ),
    .I2(\u_cpu.rf_ram.memory[30][0] ),
    .I3(\u_cpu.rf_ram.memory[31][0] ),
    .S0(_01572_),
    .S1(_01574_),
    .Z(_01584_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05093_ (.A1(_01570_),
    .A2(_01584_),
    .ZN(_01585_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05094_ (.I0(\u_cpu.rf_ram.memory[24][0] ),
    .I1(\u_cpu.rf_ram.memory[25][0] ),
    .I2(\u_cpu.rf_ram.memory[26][0] ),
    .I3(\u_cpu.rf_ram.memory[27][0] ),
    .S0(_01578_),
    .S1(_01580_),
    .Z(_01586_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05095_ (.A1(_01542_),
    .A2(_01586_),
    .B(_01418_),
    .ZN(_01587_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _05096_ (.A1(_01576_),
    .A2(_01583_),
    .B1(_01585_),
    .B2(_01587_),
    .C(_01426_),
    .ZN(_01588_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05097_ (.I(_01397_),
    .Z(_01589_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05098_ (.I(_01544_),
    .Z(_01590_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05099_ (.I(_01548_),
    .Z(_01591_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05100_ (.I0(\u_cpu.rf_ram.memory[52][0] ),
    .I1(\u_cpu.rf_ram.memory[53][0] ),
    .I2(\u_cpu.rf_ram.memory[54][0] ),
    .I3(\u_cpu.rf_ram.memory[55][0] ),
    .S0(_01590_),
    .S1(_01591_),
    .Z(_01592_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05101_ (.A1(_01589_),
    .A2(_01592_),
    .ZN(_01593_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05102_ (.I(_01540_),
    .Z(_01594_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05103_ (.I0(\u_cpu.rf_ram.memory[48][0] ),
    .I1(\u_cpu.rf_ram.memory[49][0] ),
    .I2(\u_cpu.rf_ram.memory[50][0] ),
    .I3(\u_cpu.rf_ram.memory[51][0] ),
    .S0(_01544_),
    .S1(_01548_),
    .Z(_01595_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05104_ (.A1(_01594_),
    .A2(_01595_),
    .B(_01564_),
    .ZN(_01596_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05105_ (.I(_01397_),
    .Z(_01597_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05106_ (.I(_01544_),
    .Z(_01598_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05107_ (.I0(\u_cpu.rf_ram.memory[60][0] ),
    .I1(\u_cpu.rf_ram.memory[61][0] ),
    .I2(\u_cpu.rf_ram.memory[62][0] ),
    .I3(\u_cpu.rf_ram.memory[63][0] ),
    .S0(_01598_),
    .S1(_01573_),
    .Z(_01599_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05108_ (.A1(_01597_),
    .A2(_01599_),
    .ZN(_01600_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05109_ (.I(_01540_),
    .Z(_01601_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05110_ (.I(_01543_),
    .Z(_01602_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05111_ (.I(_01547_),
    .Z(_01603_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05112_ (.I0(\u_cpu.rf_ram.memory[56][0] ),
    .I1(\u_cpu.rf_ram.memory[57][0] ),
    .I2(\u_cpu.rf_ram.memory[58][0] ),
    .I3(\u_cpu.rf_ram.memory[59][0] ),
    .S0(_01602_),
    .S1(_01603_),
    .Z(_01604_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05113_ (.I(_01416_),
    .Z(_01605_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05114_ (.A1(_01601_),
    .A2(_01604_),
    .B(_01605_),
    .ZN(_01606_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05115_ (.I(_01425_),
    .Z(_01607_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _05116_ (.A1(_01593_),
    .A2(_01596_),
    .B1(_01600_),
    .B2(_01606_),
    .C(_01607_),
    .ZN(_01608_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05117_ (.I(_01540_),
    .Z(_01609_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05118_ (.I(_01544_),
    .Z(_01610_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05119_ (.I(_01548_),
    .Z(_01611_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05120_ (.I0(\u_cpu.rf_ram.memory[40][0] ),
    .I1(\u_cpu.rf_ram.memory[41][0] ),
    .I2(\u_cpu.rf_ram.memory[42][0] ),
    .I3(\u_cpu.rf_ram.memory[43][0] ),
    .S0(_01610_),
    .S1(_01611_),
    .Z(_01612_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05121_ (.A1(_01609_),
    .A2(_01612_),
    .ZN(_01613_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05122_ (.I(_01397_),
    .Z(_01614_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05123_ (.I(_01543_),
    .Z(_01615_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05124_ (.I(_01547_),
    .Z(_01616_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05125_ (.I0(\u_cpu.rf_ram.memory[44][0] ),
    .I1(\u_cpu.rf_ram.memory[45][0] ),
    .I2(\u_cpu.rf_ram.memory[46][0] ),
    .I3(\u_cpu.rf_ram.memory[47][0] ),
    .S0(_01615_),
    .S1(_01616_),
    .Z(_01617_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05126_ (.A1(_01614_),
    .A2(_01617_),
    .B(_01605_),
    .ZN(_01618_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05127_ (.I(_01544_),
    .Z(_01619_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05128_ (.I(_01548_),
    .Z(_01620_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05129_ (.I0(\u_cpu.rf_ram.memory[36][0] ),
    .I1(\u_cpu.rf_ram.memory[37][0] ),
    .I2(\u_cpu.rf_ram.memory[38][0] ),
    .I3(\u_cpu.rf_ram.memory[39][0] ),
    .S0(_01619_),
    .S1(_01620_),
    .Z(_01621_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05130_ (.A1(_01589_),
    .A2(_01621_),
    .ZN(_01622_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05131_ (.I(_01544_),
    .Z(_01623_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05132_ (.I(_01547_),
    .Z(_01624_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05133_ (.I0(\u_cpu.rf_ram.memory[32][0] ),
    .I1(\u_cpu.rf_ram.memory[33][0] ),
    .I2(\u_cpu.rf_ram.memory[34][0] ),
    .I3(\u_cpu.rf_ram.memory[35][0] ),
    .S0(_01623_),
    .S1(_01624_),
    .Z(_01625_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05134_ (.I(_01564_),
    .Z(_01626_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05135_ (.A1(_01541_),
    .A2(_01625_),
    .B(_01626_),
    .ZN(_01627_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05136_ (.I(_01567_),
    .Z(_01628_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _05137_ (.A1(_01613_),
    .A2(_01618_),
    .B1(_01622_),
    .B2(_01627_),
    .C(_01628_),
    .ZN(_01629_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _05138_ (.A1(_01422_),
    .A2(_01608_),
    .A3(_01629_),
    .Z(_01630_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _05139_ (.A1(_01539_),
    .A2(_01569_),
    .A3(_01588_),
    .B(_01630_),
    .ZN(_01631_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05140_ (.I0(\u_cpu.rf_ram.memory[108][0] ),
    .I1(\u_cpu.rf_ram.memory[109][0] ),
    .I2(\u_cpu.rf_ram.memory[110][0] ),
    .I3(\u_cpu.rf_ram.memory[111][0] ),
    .S0(_01619_),
    .S1(_01620_),
    .Z(_01632_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05141_ (.A1(_01597_),
    .A2(_01632_),
    .ZN(_01633_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05142_ (.I0(\u_cpu.rf_ram.memory[104][0] ),
    .I1(\u_cpu.rf_ram.memory[105][0] ),
    .I2(\u_cpu.rf_ram.memory[106][0] ),
    .I3(\u_cpu.rf_ram.memory[107][0] ),
    .S0(_01615_),
    .S1(_01616_),
    .Z(_01634_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05143_ (.A1(_01594_),
    .A2(_01634_),
    .B(_01416_),
    .ZN(_01635_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05144_ (.I(_01397_),
    .Z(_01636_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05145_ (.I0(\u_cpu.rf_ram.memory[100][0] ),
    .I1(\u_cpu.rf_ram.memory[101][0] ),
    .I2(\u_cpu.rf_ram.memory[102][0] ),
    .I3(\u_cpu.rf_ram.memory[103][0] ),
    .S0(_01598_),
    .S1(_01573_),
    .Z(_01637_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05146_ (.A1(_01636_),
    .A2(_01637_),
    .ZN(_01638_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05147_ (.I0(\u_cpu.rf_ram.memory[96][0] ),
    .I1(\u_cpu.rf_ram.memory[97][0] ),
    .I2(\u_cpu.rf_ram.memory[98][0] ),
    .I3(\u_cpu.rf_ram.memory[99][0] ),
    .S0(_01602_),
    .S1(_01579_),
    .Z(_01639_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05148_ (.A1(_01601_),
    .A2(_01639_),
    .B(_01626_),
    .ZN(_01640_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _05149_ (.A1(_01633_),
    .A2(_01635_),
    .B1(_01638_),
    .B2(_01640_),
    .C(_01628_),
    .ZN(_01641_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05150_ (.I(_01548_),
    .Z(_01642_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05151_ (.I0(\u_cpu.rf_ram.memory[124][0] ),
    .I1(\u_cpu.rf_ram.memory[125][0] ),
    .I2(\u_cpu.rf_ram.memory[126][0] ),
    .I3(\u_cpu.rf_ram.memory[127][0] ),
    .S0(_01545_),
    .S1(_01642_),
    .Z(_01643_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05152_ (.A1(_01398_),
    .A2(_01643_),
    .ZN(_01644_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05153_ (.I(_01540_),
    .Z(_01645_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05154_ (.I(_01544_),
    .Z(_01646_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05155_ (.I0(\u_cpu.rf_ram.memory[120][0] ),
    .I1(\u_cpu.rf_ram.memory[121][0] ),
    .I2(\u_cpu.rf_ram.memory[122][0] ),
    .I3(\u_cpu.rf_ram.memory[123][0] ),
    .S0(_01646_),
    .S1(_01603_),
    .Z(_01647_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05156_ (.I(_01416_),
    .Z(_01648_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05157_ (.A1(_01645_),
    .A2(_01647_),
    .B(_01648_),
    .ZN(_01649_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05158_ (.I0(\u_cpu.rf_ram.memory[112][0] ),
    .I1(\u_cpu.rf_ram.memory[113][0] ),
    .I2(\u_cpu.rf_ram.memory[114][0] ),
    .I3(\u_cpu.rf_ram.memory[115][0] ),
    .S0(_01590_),
    .S1(_01591_),
    .Z(_01650_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05159_ (.A1(_01541_),
    .A2(_01650_),
    .ZN(_01651_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05160_ (.I(_01547_),
    .Z(_01652_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05161_ (.I0(\u_cpu.rf_ram.memory[116][0] ),
    .I1(\u_cpu.rf_ram.memory[117][0] ),
    .I2(\u_cpu.rf_ram.memory[118][0] ),
    .I3(\u_cpu.rf_ram.memory[119][0] ),
    .S0(_01623_),
    .S1(_01652_),
    .Z(_01653_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05162_ (.I(_01564_),
    .Z(_01654_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05163_ (.A1(_01614_),
    .A2(_01653_),
    .B(_01654_),
    .ZN(_01655_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _05164_ (.A1(_01644_),
    .A2(_01649_),
    .B1(_01651_),
    .B2(_01655_),
    .C(_01607_),
    .ZN(_01656_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _05165_ (.A1(_01422_),
    .A2(_01641_),
    .A3(_01656_),
    .ZN(_01657_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05166_ (.I0(\u_cpu.rf_ram.memory[92][0] ),
    .I1(\u_cpu.rf_ram.memory[93][0] ),
    .I2(\u_cpu.rf_ram.memory[94][0] ),
    .I3(\u_cpu.rf_ram.memory[95][0] ),
    .S0(_01610_),
    .S1(_01611_),
    .Z(_01658_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05167_ (.A1(_01398_),
    .A2(_01658_),
    .ZN(_01659_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05168_ (.I0(\u_cpu.rf_ram.memory[88][0] ),
    .I1(\u_cpu.rf_ram.memory[89][0] ),
    .I2(\u_cpu.rf_ram.memory[90][0] ),
    .I3(\u_cpu.rf_ram.memory[91][0] ),
    .S0(_01646_),
    .S1(_01624_),
    .Z(_01660_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05169_ (.A1(_01645_),
    .A2(_01660_),
    .B(_01648_),
    .ZN(_01661_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05170_ (.I0(\u_cpu.rf_ram.memory[80][0] ),
    .I1(\u_cpu.rf_ram.memory[81][0] ),
    .I2(\u_cpu.rf_ram.memory[82][0] ),
    .I3(\u_cpu.rf_ram.memory[83][0] ),
    .S0(_01545_),
    .S1(_01642_),
    .Z(_01662_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05171_ (.A1(_01609_),
    .A2(_01662_),
    .ZN(_01663_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05172_ (.I0(\u_cpu.rf_ram.memory[84][0] ),
    .I1(\u_cpu.rf_ram.memory[85][0] ),
    .I2(\u_cpu.rf_ram.memory[86][0] ),
    .I3(\u_cpu.rf_ram.memory[87][0] ),
    .S0(_01555_),
    .S1(_01652_),
    .Z(_01664_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05173_ (.A1(_01553_),
    .A2(_01664_),
    .B(_01654_),
    .ZN(_01665_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _05174_ (.A1(_01659_),
    .A2(_01661_),
    .B1(_01663_),
    .B2(_01665_),
    .C(_01426_),
    .ZN(_01666_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05175_ (.I(_01540_),
    .Z(_01667_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05176_ (.I(_01548_),
    .Z(_01668_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05177_ (.I0(\u_cpu.rf_ram.memory[64][0] ),
    .I1(\u_cpu.rf_ram.memory[65][0] ),
    .I2(\u_cpu.rf_ram.memory[66][0] ),
    .I3(\u_cpu.rf_ram.memory[67][0] ),
    .S0(_01571_),
    .S1(_01668_),
    .Z(_01669_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05178_ (.A1(_01667_),
    .A2(_01669_),
    .ZN(_01670_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05179_ (.I0(\u_cpu.rf_ram.memory[68][0] ),
    .I1(\u_cpu.rf_ram.memory[69][0] ),
    .I2(\u_cpu.rf_ram.memory[70][0] ),
    .I3(\u_cpu.rf_ram.memory[71][0] ),
    .S0(_01577_),
    .S1(_01549_),
    .Z(_01671_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05180_ (.A1(_01553_),
    .A2(_01671_),
    .B(_01565_),
    .ZN(_01672_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05181_ (.I0(\u_cpu.rf_ram.memory[72][0] ),
    .I1(\u_cpu.rf_ram.memory[73][0] ),
    .I2(\u_cpu.rf_ram.memory[74][0] ),
    .I3(\u_cpu.rf_ram.memory[75][0] ),
    .S0(_01571_),
    .S1(_01668_),
    .Z(_01673_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05182_ (.A1(_01667_),
    .A2(_01673_),
    .ZN(_01674_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05183_ (.I0(\u_cpu.rf_ram.memory[76][0] ),
    .I1(\u_cpu.rf_ram.memory[77][0] ),
    .I2(\u_cpu.rf_ram.memory[78][0] ),
    .I3(\u_cpu.rf_ram.memory[79][0] ),
    .S0(_01577_),
    .S1(_01549_),
    .Z(_01675_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05184_ (.A1(_01636_),
    .A2(_01675_),
    .B(_01417_),
    .ZN(_01676_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _05185_ (.A1(_01670_),
    .A2(_01672_),
    .B1(_01674_),
    .B2(_01676_),
    .C(_01568_),
    .ZN(_01677_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _05186_ (.A1(_01539_),
    .A2(_01666_),
    .A3(_01677_),
    .ZN(_01678_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05187_ (.A1(_01657_),
    .A2(_01678_),
    .B(_01402_),
    .ZN(_01679_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05188_ (.I(_01571_),
    .Z(_01680_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05189_ (.I(_01668_),
    .Z(_01681_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05190_ (.I0(\u_cpu.rf_ram.memory[136][0] ),
    .I1(\u_cpu.rf_ram.memory[137][0] ),
    .I2(\u_cpu.rf_ram.memory[138][0] ),
    .I3(\u_cpu.rf_ram.memory[139][0] ),
    .S0(_01680_),
    .S1(_01681_),
    .Z(_01682_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05191_ (.A1(_01399_),
    .A2(_01682_),
    .ZN(_01683_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05192_ (.I(_01667_),
    .Z(_01684_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05193_ (.I0(\u_cpu.rf_ram.memory[140][0] ),
    .I1(\u_cpu.rf_ram.memory[141][0] ),
    .I2(\u_cpu.rf_ram.memory[142][0] ),
    .I3(\u_cpu.rf_ram.memory[143][0] ),
    .S0(_01680_),
    .S1(_01681_),
    .Z(_01685_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05194_ (.A1(_01684_),
    .A2(_01685_),
    .B(_01582_),
    .ZN(_01686_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05195_ (.I(_01571_),
    .Z(_01687_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05196_ (.I(_01668_),
    .Z(_01688_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05197_ (.I0(\u_cpu.rf_ram.memory[128][0] ),
    .I1(\u_cpu.rf_ram.memory[129][0] ),
    .I2(\u_cpu.rf_ram.memory[130][0] ),
    .I3(\u_cpu.rf_ram.memory[131][0] ),
    .S0(_01687_),
    .S1(_01688_),
    .Z(_01689_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05198_ (.A1(_01399_),
    .A2(_01689_),
    .ZN(_01690_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05199_ (.I0(\u_cpu.rf_ram.memory[132][0] ),
    .I1(\u_cpu.rf_ram.memory[133][0] ),
    .I2(\u_cpu.rf_ram.memory[134][0] ),
    .I3(\u_cpu.rf_ram.memory[135][0] ),
    .S0(_01687_),
    .S1(_01688_),
    .Z(_01691_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05200_ (.A1(_01684_),
    .A2(_01691_),
    .B(_01418_),
    .ZN(_01692_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _05201_ (.A1(_01683_),
    .A2(_01686_),
    .B1(_01690_),
    .B2(_01692_),
    .C(_01404_),
    .ZN(_01693_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05202_ (.A1(_01679_),
    .A2(_01693_),
    .ZN(_01694_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05203_ (.A1(_01406_),
    .A2(_01631_),
    .B(_01694_),
    .ZN(_00000_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05204_ (.I0(\u_cpu.rf_ram.memory[8][1] ),
    .I1(\u_cpu.rf_ram.memory[9][1] ),
    .I2(\u_cpu.rf_ram.memory[10][1] ),
    .I3(\u_cpu.rf_ram.memory[11][1] ),
    .S0(_01546_),
    .S1(_01550_),
    .Z(_01695_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05205_ (.A1(_01542_),
    .A2(_01695_),
    .ZN(_01696_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05206_ (.I0(\u_cpu.rf_ram.memory[12][1] ),
    .I1(\u_cpu.rf_ram.memory[13][1] ),
    .I2(\u_cpu.rf_ram.memory[14][1] ),
    .I3(\u_cpu.rf_ram.memory[15][1] ),
    .S0(_01556_),
    .S1(_01557_),
    .Z(_01697_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05207_ (.A1(_01554_),
    .A2(_01697_),
    .B(_01417_),
    .ZN(_01698_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05208_ (.I0(\u_cpu.rf_ram.memory[4][1] ),
    .I1(\u_cpu.rf_ram.memory[5][1] ),
    .I2(\u_cpu.rf_ram.memory[6][1] ),
    .I3(\u_cpu.rf_ram.memory[7][1] ),
    .S0(_01546_),
    .S1(_01550_),
    .Z(_01699_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05209_ (.A1(_01554_),
    .A2(_01699_),
    .ZN(_01700_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05210_ (.I0(\u_cpu.rf_ram.memory[0][1] ),
    .I1(\u_cpu.rf_ram.memory[1][1] ),
    .I2(\u_cpu.rf_ram.memory[2][1] ),
    .I3(\u_cpu.rf_ram.memory[3][1] ),
    .S0(_01556_),
    .S1(_01557_),
    .Z(_01701_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05211_ (.A1(_01562_),
    .A2(_01701_),
    .B(_01565_),
    .ZN(_01702_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _05212_ (.A1(_01696_),
    .A2(_01698_),
    .B1(_01700_),
    .B2(_01702_),
    .C(_01568_),
    .ZN(_01703_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05213_ (.I0(\u_cpu.rf_ram.memory[20][1] ),
    .I1(\u_cpu.rf_ram.memory[21][1] ),
    .I2(\u_cpu.rf_ram.memory[22][1] ),
    .I3(\u_cpu.rf_ram.memory[23][1] ),
    .S0(_01572_),
    .S1(_01574_),
    .Z(_01704_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05214_ (.A1(_01570_),
    .A2(_01704_),
    .ZN(_01705_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05215_ (.I0(\u_cpu.rf_ram.memory[16][1] ),
    .I1(\u_cpu.rf_ram.memory[17][1] ),
    .I2(\u_cpu.rf_ram.memory[18][1] ),
    .I3(\u_cpu.rf_ram.memory[19][1] ),
    .S0(_01578_),
    .S1(_01580_),
    .Z(_01706_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05216_ (.A1(_01562_),
    .A2(_01706_),
    .B(_01582_),
    .ZN(_01707_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05217_ (.I0(\u_cpu.rf_ram.memory[28][1] ),
    .I1(\u_cpu.rf_ram.memory[29][1] ),
    .I2(\u_cpu.rf_ram.memory[30][1] ),
    .I3(\u_cpu.rf_ram.memory[31][1] ),
    .S0(_01572_),
    .S1(_01574_),
    .Z(_01708_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05218_ (.A1(_01570_),
    .A2(_01708_),
    .ZN(_01709_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05219_ (.I0(\u_cpu.rf_ram.memory[24][1] ),
    .I1(\u_cpu.rf_ram.memory[25][1] ),
    .I2(\u_cpu.rf_ram.memory[26][1] ),
    .I3(\u_cpu.rf_ram.memory[27][1] ),
    .S0(_01578_),
    .S1(_01580_),
    .Z(_01710_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05220_ (.A1(_01542_),
    .A2(_01710_),
    .B(_01418_),
    .ZN(_01711_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _05221_ (.A1(_01705_),
    .A2(_01707_),
    .B1(_01709_),
    .B2(_01711_),
    .C(_01426_),
    .ZN(_01712_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05222_ (.I0(\u_cpu.rf_ram.memory[52][1] ),
    .I1(\u_cpu.rf_ram.memory[53][1] ),
    .I2(\u_cpu.rf_ram.memory[54][1] ),
    .I3(\u_cpu.rf_ram.memory[55][1] ),
    .S0(_01590_),
    .S1(_01591_),
    .Z(_01713_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05223_ (.A1(_01589_),
    .A2(_01713_),
    .ZN(_01714_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05224_ (.I0(\u_cpu.rf_ram.memory[48][1] ),
    .I1(\u_cpu.rf_ram.memory[49][1] ),
    .I2(\u_cpu.rf_ram.memory[50][1] ),
    .I3(\u_cpu.rf_ram.memory[51][1] ),
    .S0(_01544_),
    .S1(_01548_),
    .Z(_01715_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05225_ (.A1(_01594_),
    .A2(_01715_),
    .B(_01564_),
    .ZN(_01716_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05226_ (.I0(\u_cpu.rf_ram.memory[60][1] ),
    .I1(\u_cpu.rf_ram.memory[61][1] ),
    .I2(\u_cpu.rf_ram.memory[62][1] ),
    .I3(\u_cpu.rf_ram.memory[63][1] ),
    .S0(_01598_),
    .S1(_01573_),
    .Z(_01717_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05227_ (.A1(_01597_),
    .A2(_01717_),
    .ZN(_01718_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05228_ (.I0(\u_cpu.rf_ram.memory[56][1] ),
    .I1(\u_cpu.rf_ram.memory[57][1] ),
    .I2(\u_cpu.rf_ram.memory[58][1] ),
    .I3(\u_cpu.rf_ram.memory[59][1] ),
    .S0(_01602_),
    .S1(_01579_),
    .Z(_01719_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05229_ (.A1(_01601_),
    .A2(_01719_),
    .B(_01605_),
    .ZN(_01720_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _05230_ (.A1(_01714_),
    .A2(_01716_),
    .B1(_01718_),
    .B2(_01720_),
    .C(_01607_),
    .ZN(_01721_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05231_ (.I0(\u_cpu.rf_ram.memory[40][1] ),
    .I1(\u_cpu.rf_ram.memory[41][1] ),
    .I2(\u_cpu.rf_ram.memory[42][1] ),
    .I3(\u_cpu.rf_ram.memory[43][1] ),
    .S0(_01610_),
    .S1(_01611_),
    .Z(_01722_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05232_ (.A1(_01609_),
    .A2(_01722_),
    .ZN(_01723_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05233_ (.I0(\u_cpu.rf_ram.memory[44][1] ),
    .I1(\u_cpu.rf_ram.memory[45][1] ),
    .I2(\u_cpu.rf_ram.memory[46][1] ),
    .I3(\u_cpu.rf_ram.memory[47][1] ),
    .S0(_01615_),
    .S1(_01616_),
    .Z(_01724_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05234_ (.A1(_01614_),
    .A2(_01724_),
    .B(_01605_),
    .ZN(_01725_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05235_ (.I0(\u_cpu.rf_ram.memory[36][1] ),
    .I1(\u_cpu.rf_ram.memory[37][1] ),
    .I2(\u_cpu.rf_ram.memory[38][1] ),
    .I3(\u_cpu.rf_ram.memory[39][1] ),
    .S0(_01619_),
    .S1(_01620_),
    .Z(_01726_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05236_ (.A1(_01589_),
    .A2(_01726_),
    .ZN(_01727_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05237_ (.I0(\u_cpu.rf_ram.memory[32][1] ),
    .I1(\u_cpu.rf_ram.memory[33][1] ),
    .I2(\u_cpu.rf_ram.memory[34][1] ),
    .I3(\u_cpu.rf_ram.memory[35][1] ),
    .S0(_01623_),
    .S1(_01624_),
    .Z(_01728_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05238_ (.A1(_01541_),
    .A2(_01728_),
    .B(_01626_),
    .ZN(_01729_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _05239_ (.A1(_01723_),
    .A2(_01725_),
    .B1(_01727_),
    .B2(_01729_),
    .C(_01628_),
    .ZN(_01730_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _05240_ (.A1(_01422_),
    .A2(_01721_),
    .A3(_01730_),
    .Z(_01731_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _05241_ (.A1(_01539_),
    .A2(_01703_),
    .A3(_01712_),
    .B(_01731_),
    .ZN(_01732_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05242_ (.I0(\u_cpu.rf_ram.memory[108][1] ),
    .I1(\u_cpu.rf_ram.memory[109][1] ),
    .I2(\u_cpu.rf_ram.memory[110][1] ),
    .I3(\u_cpu.rf_ram.memory[111][1] ),
    .S0(_01619_),
    .S1(_01620_),
    .Z(_01733_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05243_ (.A1(_01597_),
    .A2(_01733_),
    .ZN(_01734_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05244_ (.I0(\u_cpu.rf_ram.memory[104][1] ),
    .I1(\u_cpu.rf_ram.memory[105][1] ),
    .I2(\u_cpu.rf_ram.memory[106][1] ),
    .I3(\u_cpu.rf_ram.memory[107][1] ),
    .S0(_01615_),
    .S1(_01616_),
    .Z(_01735_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05245_ (.A1(_01594_),
    .A2(_01735_),
    .B(_01416_),
    .ZN(_01736_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05246_ (.I0(\u_cpu.rf_ram.memory[100][1] ),
    .I1(\u_cpu.rf_ram.memory[101][1] ),
    .I2(\u_cpu.rf_ram.memory[102][1] ),
    .I3(\u_cpu.rf_ram.memory[103][1] ),
    .S0(_01598_),
    .S1(_01573_),
    .Z(_01737_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05247_ (.A1(_01636_),
    .A2(_01737_),
    .ZN(_01738_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05248_ (.I0(\u_cpu.rf_ram.memory[96][1] ),
    .I1(\u_cpu.rf_ram.memory[97][1] ),
    .I2(\u_cpu.rf_ram.memory[98][1] ),
    .I3(\u_cpu.rf_ram.memory[99][1] ),
    .S0(_01602_),
    .S1(_01579_),
    .Z(_01739_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05249_ (.A1(_01601_),
    .A2(_01739_),
    .B(_01626_),
    .ZN(_01740_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _05250_ (.A1(_01734_),
    .A2(_01736_),
    .B1(_01738_),
    .B2(_01740_),
    .C(_01628_),
    .ZN(_01741_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05251_ (.I0(\u_cpu.rf_ram.memory[124][1] ),
    .I1(\u_cpu.rf_ram.memory[125][1] ),
    .I2(\u_cpu.rf_ram.memory[126][1] ),
    .I3(\u_cpu.rf_ram.memory[127][1] ),
    .S0(_01545_),
    .S1(_01642_),
    .Z(_01742_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05252_ (.A1(_01398_),
    .A2(_01742_),
    .ZN(_01743_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05253_ (.I0(\u_cpu.rf_ram.memory[120][1] ),
    .I1(\u_cpu.rf_ram.memory[121][1] ),
    .I2(\u_cpu.rf_ram.memory[122][1] ),
    .I3(\u_cpu.rf_ram.memory[123][1] ),
    .S0(_01646_),
    .S1(_01603_),
    .Z(_01744_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05254_ (.A1(_01645_),
    .A2(_01744_),
    .B(_01648_),
    .ZN(_01745_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05255_ (.I0(\u_cpu.rf_ram.memory[112][1] ),
    .I1(\u_cpu.rf_ram.memory[113][1] ),
    .I2(\u_cpu.rf_ram.memory[114][1] ),
    .I3(\u_cpu.rf_ram.memory[115][1] ),
    .S0(_01590_),
    .S1(_01591_),
    .Z(_01746_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05256_ (.A1(_01541_),
    .A2(_01746_),
    .ZN(_01747_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05257_ (.I0(\u_cpu.rf_ram.memory[116][1] ),
    .I1(\u_cpu.rf_ram.memory[117][1] ),
    .I2(\u_cpu.rf_ram.memory[118][1] ),
    .I3(\u_cpu.rf_ram.memory[119][1] ),
    .S0(_01623_),
    .S1(_01624_),
    .Z(_01748_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05258_ (.A1(_01614_),
    .A2(_01748_),
    .B(_01654_),
    .ZN(_01749_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _05259_ (.A1(_01743_),
    .A2(_01745_),
    .B1(_01747_),
    .B2(_01749_),
    .C(_01607_),
    .ZN(_01750_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _05260_ (.A1(_01422_),
    .A2(_01741_),
    .A3(_01750_),
    .ZN(_01751_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05261_ (.I0(\u_cpu.rf_ram.memory[92][1] ),
    .I1(\u_cpu.rf_ram.memory[93][1] ),
    .I2(\u_cpu.rf_ram.memory[94][1] ),
    .I3(\u_cpu.rf_ram.memory[95][1] ),
    .S0(_01610_),
    .S1(_01611_),
    .Z(_01752_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05262_ (.A1(_01398_),
    .A2(_01752_),
    .ZN(_01753_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05263_ (.I0(\u_cpu.rf_ram.memory[88][1] ),
    .I1(\u_cpu.rf_ram.memory[89][1] ),
    .I2(\u_cpu.rf_ram.memory[90][1] ),
    .I3(\u_cpu.rf_ram.memory[91][1] ),
    .S0(_01646_),
    .S1(_01603_),
    .Z(_01754_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05264_ (.A1(_01645_),
    .A2(_01754_),
    .B(_01648_),
    .ZN(_01755_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05265_ (.I0(\u_cpu.rf_ram.memory[80][1] ),
    .I1(\u_cpu.rf_ram.memory[81][1] ),
    .I2(\u_cpu.rf_ram.memory[82][1] ),
    .I3(\u_cpu.rf_ram.memory[83][1] ),
    .S0(_01545_),
    .S1(_01642_),
    .Z(_01756_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05266_ (.A1(_01609_),
    .A2(_01756_),
    .ZN(_01757_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05267_ (.I0(\u_cpu.rf_ram.memory[84][1] ),
    .I1(\u_cpu.rf_ram.memory[85][1] ),
    .I2(\u_cpu.rf_ram.memory[86][1] ),
    .I3(\u_cpu.rf_ram.memory[87][1] ),
    .S0(_01555_),
    .S1(_01652_),
    .Z(_01758_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05268_ (.A1(_01553_),
    .A2(_01758_),
    .B(_01654_),
    .ZN(_01759_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _05269_ (.A1(_01753_),
    .A2(_01755_),
    .B1(_01757_),
    .B2(_01759_),
    .C(_01426_),
    .ZN(_01760_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05270_ (.I0(\u_cpu.rf_ram.memory[64][1] ),
    .I1(\u_cpu.rf_ram.memory[65][1] ),
    .I2(\u_cpu.rf_ram.memory[66][1] ),
    .I3(\u_cpu.rf_ram.memory[67][1] ),
    .S0(_01571_),
    .S1(_01668_),
    .Z(_01761_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05271_ (.A1(_01667_),
    .A2(_01761_),
    .ZN(_01762_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05272_ (.I0(\u_cpu.rf_ram.memory[68][1] ),
    .I1(\u_cpu.rf_ram.memory[69][1] ),
    .I2(\u_cpu.rf_ram.memory[70][1] ),
    .I3(\u_cpu.rf_ram.memory[71][1] ),
    .S0(_01555_),
    .S1(_01652_),
    .Z(_01763_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05273_ (.A1(_01553_),
    .A2(_01763_),
    .B(_01565_),
    .ZN(_01764_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05274_ (.I0(\u_cpu.rf_ram.memory[72][1] ),
    .I1(\u_cpu.rf_ram.memory[73][1] ),
    .I2(\u_cpu.rf_ram.memory[74][1] ),
    .I3(\u_cpu.rf_ram.memory[75][1] ),
    .S0(_01571_),
    .S1(_01668_),
    .Z(_01765_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05275_ (.A1(_01667_),
    .A2(_01765_),
    .ZN(_01766_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05276_ (.I0(\u_cpu.rf_ram.memory[76][1] ),
    .I1(\u_cpu.rf_ram.memory[77][1] ),
    .I2(\u_cpu.rf_ram.memory[78][1] ),
    .I3(\u_cpu.rf_ram.memory[79][1] ),
    .S0(_01577_),
    .S1(_01549_),
    .Z(_01767_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05277_ (.A1(_01636_),
    .A2(_01767_),
    .B(_01417_),
    .ZN(_01768_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _05278_ (.A1(_01762_),
    .A2(_01764_),
    .B1(_01766_),
    .B2(_01768_),
    .C(_01568_),
    .ZN(_01769_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _05279_ (.A1(_01539_),
    .A2(_01760_),
    .A3(_01769_),
    .ZN(_01770_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05280_ (.A1(_01751_),
    .A2(_01770_),
    .B(_01402_),
    .ZN(_01771_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05281_ (.I0(\u_cpu.rf_ram.memory[136][1] ),
    .I1(\u_cpu.rf_ram.memory[137][1] ),
    .I2(\u_cpu.rf_ram.memory[138][1] ),
    .I3(\u_cpu.rf_ram.memory[139][1] ),
    .S0(_01680_),
    .S1(_01681_),
    .Z(_01772_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05282_ (.A1(_01399_),
    .A2(_01772_),
    .ZN(_01773_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05283_ (.I0(\u_cpu.rf_ram.memory[140][1] ),
    .I1(\u_cpu.rf_ram.memory[141][1] ),
    .I2(\u_cpu.rf_ram.memory[142][1] ),
    .I3(\u_cpu.rf_ram.memory[143][1] ),
    .S0(_01680_),
    .S1(_01681_),
    .Z(_01774_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05284_ (.A1(_01684_),
    .A2(_01774_),
    .B(_01582_),
    .ZN(_01775_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05285_ (.I0(\u_cpu.rf_ram.memory[128][1] ),
    .I1(\u_cpu.rf_ram.memory[129][1] ),
    .I2(\u_cpu.rf_ram.memory[130][1] ),
    .I3(\u_cpu.rf_ram.memory[131][1] ),
    .S0(_01687_),
    .S1(_01688_),
    .Z(_01776_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05286_ (.A1(_01399_),
    .A2(_01776_),
    .ZN(_01777_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05287_ (.I0(\u_cpu.rf_ram.memory[132][1] ),
    .I1(\u_cpu.rf_ram.memory[133][1] ),
    .I2(\u_cpu.rf_ram.memory[134][1] ),
    .I3(\u_cpu.rf_ram.memory[135][1] ),
    .S0(_01687_),
    .S1(_01688_),
    .Z(_01778_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05288_ (.A1(_01684_),
    .A2(_01778_),
    .B(_01418_),
    .ZN(_01779_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _05289_ (.A1(_01773_),
    .A2(_01775_),
    .B1(_01777_),
    .B2(_01779_),
    .C(_01404_),
    .ZN(_01780_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05290_ (.A1(_01771_),
    .A2(_01780_),
    .ZN(_01781_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05291_ (.A1(_01406_),
    .A2(_01732_),
    .B(_01781_),
    .ZN(_00001_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05292_ (.I0(\u_cpu.rf_ram.memory[8][2] ),
    .I1(\u_cpu.rf_ram.memory[9][2] ),
    .I2(\u_cpu.rf_ram.memory[10][2] ),
    .I3(\u_cpu.rf_ram.memory[11][2] ),
    .S0(_01546_),
    .S1(_01550_),
    .Z(_01782_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05293_ (.A1(_01542_),
    .A2(_01782_),
    .ZN(_01783_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05294_ (.I0(\u_cpu.rf_ram.memory[12][2] ),
    .I1(\u_cpu.rf_ram.memory[13][2] ),
    .I2(\u_cpu.rf_ram.memory[14][2] ),
    .I3(\u_cpu.rf_ram.memory[15][2] ),
    .S0(_01556_),
    .S1(_01557_),
    .Z(_01784_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05295_ (.A1(_01554_),
    .A2(_01784_),
    .B(_01417_),
    .ZN(_01785_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05296_ (.I0(\u_cpu.rf_ram.memory[4][2] ),
    .I1(\u_cpu.rf_ram.memory[5][2] ),
    .I2(\u_cpu.rf_ram.memory[6][2] ),
    .I3(\u_cpu.rf_ram.memory[7][2] ),
    .S0(_01546_),
    .S1(_01550_),
    .Z(_01786_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05297_ (.A1(_01554_),
    .A2(_01786_),
    .ZN(_01787_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05298_ (.I0(\u_cpu.rf_ram.memory[0][2] ),
    .I1(\u_cpu.rf_ram.memory[1][2] ),
    .I2(\u_cpu.rf_ram.memory[2][2] ),
    .I3(\u_cpu.rf_ram.memory[3][2] ),
    .S0(_01556_),
    .S1(_01557_),
    .Z(_01788_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05299_ (.A1(_01562_),
    .A2(_01788_),
    .B(_01565_),
    .ZN(_01789_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _05300_ (.A1(_01783_),
    .A2(_01785_),
    .B1(_01787_),
    .B2(_01789_),
    .C(_01568_),
    .ZN(_01790_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05301_ (.I0(\u_cpu.rf_ram.memory[20][2] ),
    .I1(\u_cpu.rf_ram.memory[21][2] ),
    .I2(\u_cpu.rf_ram.memory[22][2] ),
    .I3(\u_cpu.rf_ram.memory[23][2] ),
    .S0(_01572_),
    .S1(_01574_),
    .Z(_01791_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05302_ (.A1(_01570_),
    .A2(_01791_),
    .ZN(_01792_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05303_ (.I0(\u_cpu.rf_ram.memory[16][2] ),
    .I1(\u_cpu.rf_ram.memory[17][2] ),
    .I2(\u_cpu.rf_ram.memory[18][2] ),
    .I3(\u_cpu.rf_ram.memory[19][2] ),
    .S0(_01578_),
    .S1(_01580_),
    .Z(_01793_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05304_ (.A1(_01562_),
    .A2(_01793_),
    .B(_01582_),
    .ZN(_01794_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05305_ (.I0(\u_cpu.rf_ram.memory[28][2] ),
    .I1(\u_cpu.rf_ram.memory[29][2] ),
    .I2(\u_cpu.rf_ram.memory[30][2] ),
    .I3(\u_cpu.rf_ram.memory[31][2] ),
    .S0(_01572_),
    .S1(_01574_),
    .Z(_01795_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05306_ (.A1(_01570_),
    .A2(_01795_),
    .ZN(_01796_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05307_ (.I0(\u_cpu.rf_ram.memory[24][2] ),
    .I1(\u_cpu.rf_ram.memory[25][2] ),
    .I2(\u_cpu.rf_ram.memory[26][2] ),
    .I3(\u_cpu.rf_ram.memory[27][2] ),
    .S0(_01578_),
    .S1(_01580_),
    .Z(_01797_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05308_ (.A1(_01542_),
    .A2(_01797_),
    .B(_01418_),
    .ZN(_01798_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _05309_ (.A1(_01792_),
    .A2(_01794_),
    .B1(_01796_),
    .B2(_01798_),
    .C(_01426_),
    .ZN(_01799_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05310_ (.I0(\u_cpu.rf_ram.memory[52][2] ),
    .I1(\u_cpu.rf_ram.memory[53][2] ),
    .I2(\u_cpu.rf_ram.memory[54][2] ),
    .I3(\u_cpu.rf_ram.memory[55][2] ),
    .S0(_01590_),
    .S1(_01591_),
    .Z(_01800_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05311_ (.A1(_01589_),
    .A2(_01800_),
    .ZN(_01801_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05312_ (.I0(\u_cpu.rf_ram.memory[48][2] ),
    .I1(\u_cpu.rf_ram.memory[49][2] ),
    .I2(\u_cpu.rf_ram.memory[50][2] ),
    .I3(\u_cpu.rf_ram.memory[51][2] ),
    .S0(_01544_),
    .S1(_01548_),
    .Z(_01802_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05313_ (.A1(_01594_),
    .A2(_01802_),
    .B(_01564_),
    .ZN(_01803_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05314_ (.I0(\u_cpu.rf_ram.memory[60][2] ),
    .I1(\u_cpu.rf_ram.memory[61][2] ),
    .I2(\u_cpu.rf_ram.memory[62][2] ),
    .I3(\u_cpu.rf_ram.memory[63][2] ),
    .S0(_01598_),
    .S1(_01573_),
    .Z(_01804_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05315_ (.A1(_01597_),
    .A2(_01804_),
    .ZN(_01805_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05316_ (.I0(\u_cpu.rf_ram.memory[56][2] ),
    .I1(\u_cpu.rf_ram.memory[57][2] ),
    .I2(\u_cpu.rf_ram.memory[58][2] ),
    .I3(\u_cpu.rf_ram.memory[59][2] ),
    .S0(_01602_),
    .S1(_01579_),
    .Z(_01806_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05317_ (.A1(_01601_),
    .A2(_01806_),
    .B(_01605_),
    .ZN(_01807_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _05318_ (.A1(_01801_),
    .A2(_01803_),
    .B1(_01805_),
    .B2(_01807_),
    .C(_01607_),
    .ZN(_01808_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05319_ (.I0(\u_cpu.rf_ram.memory[40][2] ),
    .I1(\u_cpu.rf_ram.memory[41][2] ),
    .I2(\u_cpu.rf_ram.memory[42][2] ),
    .I3(\u_cpu.rf_ram.memory[43][2] ),
    .S0(_01610_),
    .S1(_01611_),
    .Z(_01809_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05320_ (.A1(_01609_),
    .A2(_01809_),
    .ZN(_01810_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05321_ (.I0(\u_cpu.rf_ram.memory[44][2] ),
    .I1(\u_cpu.rf_ram.memory[45][2] ),
    .I2(\u_cpu.rf_ram.memory[46][2] ),
    .I3(\u_cpu.rf_ram.memory[47][2] ),
    .S0(_01615_),
    .S1(_01616_),
    .Z(_01811_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05322_ (.A1(_01614_),
    .A2(_01811_),
    .B(_01605_),
    .ZN(_01812_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05323_ (.I0(\u_cpu.rf_ram.memory[36][2] ),
    .I1(\u_cpu.rf_ram.memory[37][2] ),
    .I2(\u_cpu.rf_ram.memory[38][2] ),
    .I3(\u_cpu.rf_ram.memory[39][2] ),
    .S0(_01619_),
    .S1(_01620_),
    .Z(_01813_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05324_ (.A1(_01589_),
    .A2(_01813_),
    .ZN(_01814_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05325_ (.I0(\u_cpu.rf_ram.memory[32][2] ),
    .I1(\u_cpu.rf_ram.memory[33][2] ),
    .I2(\u_cpu.rf_ram.memory[34][2] ),
    .I3(\u_cpu.rf_ram.memory[35][2] ),
    .S0(_01623_),
    .S1(_01624_),
    .Z(_01815_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05326_ (.A1(_01541_),
    .A2(_01815_),
    .B(_01626_),
    .ZN(_01816_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _05327_ (.A1(_01810_),
    .A2(_01812_),
    .B1(_01814_),
    .B2(_01816_),
    .C(_01628_),
    .ZN(_01817_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _05328_ (.A1(_01422_),
    .A2(_01808_),
    .A3(_01817_),
    .Z(_01818_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _05329_ (.A1(_01539_),
    .A2(_01790_),
    .A3(_01799_),
    .B(_01818_),
    .ZN(_01819_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05330_ (.I0(\u_cpu.rf_ram.memory[108][2] ),
    .I1(\u_cpu.rf_ram.memory[109][2] ),
    .I2(\u_cpu.rf_ram.memory[110][2] ),
    .I3(\u_cpu.rf_ram.memory[111][2] ),
    .S0(_01598_),
    .S1(_01620_),
    .Z(_01820_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05331_ (.A1(_01597_),
    .A2(_01820_),
    .ZN(_01821_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05332_ (.I0(\u_cpu.rf_ram.memory[104][2] ),
    .I1(\u_cpu.rf_ram.memory[105][2] ),
    .I2(\u_cpu.rf_ram.memory[106][2] ),
    .I3(\u_cpu.rf_ram.memory[107][2] ),
    .S0(_01615_),
    .S1(_01616_),
    .Z(_01822_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05333_ (.A1(_01594_),
    .A2(_01822_),
    .B(_01416_),
    .ZN(_01823_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05334_ (.I0(\u_cpu.rf_ram.memory[100][2] ),
    .I1(\u_cpu.rf_ram.memory[101][2] ),
    .I2(\u_cpu.rf_ram.memory[102][2] ),
    .I3(\u_cpu.rf_ram.memory[103][2] ),
    .S0(_01577_),
    .S1(_01549_),
    .Z(_01824_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05335_ (.A1(_01636_),
    .A2(_01824_),
    .ZN(_01825_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05336_ (.I0(\u_cpu.rf_ram.memory[96][2] ),
    .I1(\u_cpu.rf_ram.memory[97][2] ),
    .I2(\u_cpu.rf_ram.memory[98][2] ),
    .I3(\u_cpu.rf_ram.memory[99][2] ),
    .S0(_01602_),
    .S1(_01579_),
    .Z(_01826_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05337_ (.A1(_01601_),
    .A2(_01826_),
    .B(_01626_),
    .ZN(_01827_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _05338_ (.A1(_01821_),
    .A2(_01823_),
    .B1(_01825_),
    .B2(_01827_),
    .C(_01628_),
    .ZN(_01828_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05339_ (.I0(\u_cpu.rf_ram.memory[124][2] ),
    .I1(\u_cpu.rf_ram.memory[125][2] ),
    .I2(\u_cpu.rf_ram.memory[126][2] ),
    .I3(\u_cpu.rf_ram.memory[127][2] ),
    .S0(_01545_),
    .S1(_01642_),
    .Z(_01829_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05340_ (.A1(_01398_),
    .A2(_01829_),
    .ZN(_01830_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05341_ (.I0(\u_cpu.rf_ram.memory[120][2] ),
    .I1(\u_cpu.rf_ram.memory[121][2] ),
    .I2(\u_cpu.rf_ram.memory[122][2] ),
    .I3(\u_cpu.rf_ram.memory[123][2] ),
    .S0(_01646_),
    .S1(_01603_),
    .Z(_01831_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05342_ (.A1(_01645_),
    .A2(_01831_),
    .B(_01648_),
    .ZN(_01832_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05343_ (.I0(\u_cpu.rf_ram.memory[112][2] ),
    .I1(\u_cpu.rf_ram.memory[113][2] ),
    .I2(\u_cpu.rf_ram.memory[114][2] ),
    .I3(\u_cpu.rf_ram.memory[115][2] ),
    .S0(_01619_),
    .S1(_01591_),
    .Z(_01833_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05344_ (.A1(_01541_),
    .A2(_01833_),
    .ZN(_01834_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05345_ (.I0(\u_cpu.rf_ram.memory[116][2] ),
    .I1(\u_cpu.rf_ram.memory[117][2] ),
    .I2(\u_cpu.rf_ram.memory[118][2] ),
    .I3(\u_cpu.rf_ram.memory[119][2] ),
    .S0(_01623_),
    .S1(_01624_),
    .Z(_01835_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05346_ (.A1(_01614_),
    .A2(_01835_),
    .B(_01654_),
    .ZN(_01836_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _05347_ (.A1(_01830_),
    .A2(_01832_),
    .B1(_01834_),
    .B2(_01836_),
    .C(_01607_),
    .ZN(_01837_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _05348_ (.A1(_01422_),
    .A2(_01828_),
    .A3(_01837_),
    .ZN(_01838_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05349_ (.I0(\u_cpu.rf_ram.memory[92][2] ),
    .I1(\u_cpu.rf_ram.memory[93][2] ),
    .I2(\u_cpu.rf_ram.memory[94][2] ),
    .I3(\u_cpu.rf_ram.memory[95][2] ),
    .S0(_01610_),
    .S1(_01611_),
    .Z(_01839_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05350_ (.A1(_01398_),
    .A2(_01839_),
    .ZN(_01840_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05351_ (.I0(\u_cpu.rf_ram.memory[88][2] ),
    .I1(\u_cpu.rf_ram.memory[89][2] ),
    .I2(\u_cpu.rf_ram.memory[90][2] ),
    .I3(\u_cpu.rf_ram.memory[91][2] ),
    .S0(_01646_),
    .S1(_01603_),
    .Z(_01841_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05352_ (.A1(_01645_),
    .A2(_01841_),
    .B(_01648_),
    .ZN(_01842_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05353_ (.I0(\u_cpu.rf_ram.memory[80][2] ),
    .I1(\u_cpu.rf_ram.memory[81][2] ),
    .I2(\u_cpu.rf_ram.memory[82][2] ),
    .I3(\u_cpu.rf_ram.memory[83][2] ),
    .S0(_01590_),
    .S1(_01642_),
    .Z(_01843_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05354_ (.A1(_01609_),
    .A2(_01843_),
    .ZN(_01844_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05355_ (.I0(\u_cpu.rf_ram.memory[84][2] ),
    .I1(\u_cpu.rf_ram.memory[85][2] ),
    .I2(\u_cpu.rf_ram.memory[86][2] ),
    .I3(\u_cpu.rf_ram.memory[87][2] ),
    .S0(_01555_),
    .S1(_01652_),
    .Z(_01845_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05356_ (.A1(_01553_),
    .A2(_01845_),
    .B(_01654_),
    .ZN(_01846_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _05357_ (.A1(_01840_),
    .A2(_01842_),
    .B1(_01844_),
    .B2(_01846_),
    .C(_01426_),
    .ZN(_01847_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05358_ (.I0(\u_cpu.rf_ram.memory[64][2] ),
    .I1(\u_cpu.rf_ram.memory[65][2] ),
    .I2(\u_cpu.rf_ram.memory[66][2] ),
    .I3(\u_cpu.rf_ram.memory[67][2] ),
    .S0(_01571_),
    .S1(_01668_),
    .Z(_01848_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05359_ (.A1(_01667_),
    .A2(_01848_),
    .ZN(_01849_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05360_ (.I0(\u_cpu.rf_ram.memory[68][2] ),
    .I1(\u_cpu.rf_ram.memory[69][2] ),
    .I2(\u_cpu.rf_ram.memory[70][2] ),
    .I3(\u_cpu.rf_ram.memory[71][2] ),
    .S0(_01555_),
    .S1(_01652_),
    .Z(_01850_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05361_ (.A1(_01553_),
    .A2(_01850_),
    .B(_01565_),
    .ZN(_01851_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05362_ (.I0(\u_cpu.rf_ram.memory[72][2] ),
    .I1(\u_cpu.rf_ram.memory[73][2] ),
    .I2(\u_cpu.rf_ram.memory[74][2] ),
    .I3(\u_cpu.rf_ram.memory[75][2] ),
    .S0(_01571_),
    .S1(_01668_),
    .Z(_01852_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05363_ (.A1(_01667_),
    .A2(_01852_),
    .ZN(_01853_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05364_ (.I0(\u_cpu.rf_ram.memory[76][2] ),
    .I1(\u_cpu.rf_ram.memory[77][2] ),
    .I2(\u_cpu.rf_ram.memory[78][2] ),
    .I3(\u_cpu.rf_ram.memory[79][2] ),
    .S0(_01577_),
    .S1(_01549_),
    .Z(_01854_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05365_ (.A1(_01636_),
    .A2(_01854_),
    .B(_01417_),
    .ZN(_01855_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _05366_ (.A1(_01849_),
    .A2(_01851_),
    .B1(_01853_),
    .B2(_01855_),
    .C(_01568_),
    .ZN(_01856_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _05367_ (.A1(_01539_),
    .A2(_01847_),
    .A3(_01856_),
    .ZN(_01857_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05368_ (.A1(_01838_),
    .A2(_01857_),
    .B(_01402_),
    .ZN(_01858_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05369_ (.I0(\u_cpu.rf_ram.memory[136][2] ),
    .I1(\u_cpu.rf_ram.memory[137][2] ),
    .I2(\u_cpu.rf_ram.memory[138][2] ),
    .I3(\u_cpu.rf_ram.memory[139][2] ),
    .S0(_01680_),
    .S1(_01681_),
    .Z(_01859_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05370_ (.A1(_01399_),
    .A2(_01859_),
    .ZN(_01860_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05371_ (.I0(\u_cpu.rf_ram.memory[140][2] ),
    .I1(\u_cpu.rf_ram.memory[141][2] ),
    .I2(\u_cpu.rf_ram.memory[142][2] ),
    .I3(\u_cpu.rf_ram.memory[143][2] ),
    .S0(_01680_),
    .S1(_01681_),
    .Z(_01861_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05372_ (.A1(_01684_),
    .A2(_01861_),
    .B(_01582_),
    .ZN(_01862_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05373_ (.I0(\u_cpu.rf_ram.memory[128][2] ),
    .I1(\u_cpu.rf_ram.memory[129][2] ),
    .I2(\u_cpu.rf_ram.memory[130][2] ),
    .I3(\u_cpu.rf_ram.memory[131][2] ),
    .S0(_01687_),
    .S1(_01688_),
    .Z(_01863_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05374_ (.A1(_01399_),
    .A2(_01863_),
    .ZN(_01864_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05375_ (.I0(\u_cpu.rf_ram.memory[132][2] ),
    .I1(\u_cpu.rf_ram.memory[133][2] ),
    .I2(\u_cpu.rf_ram.memory[134][2] ),
    .I3(\u_cpu.rf_ram.memory[135][2] ),
    .S0(_01687_),
    .S1(_01688_),
    .Z(_01865_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05376_ (.A1(_01684_),
    .A2(_01865_),
    .B(_01418_),
    .ZN(_01866_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _05377_ (.A1(_01860_),
    .A2(_01862_),
    .B1(_01864_),
    .B2(_01866_),
    .C(_01404_),
    .ZN(_01867_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05378_ (.A1(_01858_),
    .A2(_01867_),
    .ZN(_01868_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05379_ (.A1(_01406_),
    .A2(_01819_),
    .B(_01868_),
    .ZN(_00002_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05380_ (.I0(\u_cpu.rf_ram.memory[8][3] ),
    .I1(\u_cpu.rf_ram.memory[9][3] ),
    .I2(\u_cpu.rf_ram.memory[10][3] ),
    .I3(\u_cpu.rf_ram.memory[11][3] ),
    .S0(_01546_),
    .S1(_01550_),
    .Z(_01869_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05381_ (.A1(_01542_),
    .A2(_01869_),
    .ZN(_01870_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05382_ (.I0(\u_cpu.rf_ram.memory[12][3] ),
    .I1(\u_cpu.rf_ram.memory[13][3] ),
    .I2(\u_cpu.rf_ram.memory[14][3] ),
    .I3(\u_cpu.rf_ram.memory[15][3] ),
    .S0(_01556_),
    .S1(_01557_),
    .Z(_01871_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05383_ (.A1(_01554_),
    .A2(_01871_),
    .B(_01417_),
    .ZN(_01872_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05384_ (.I0(\u_cpu.rf_ram.memory[4][3] ),
    .I1(\u_cpu.rf_ram.memory[5][3] ),
    .I2(\u_cpu.rf_ram.memory[6][3] ),
    .I3(\u_cpu.rf_ram.memory[7][3] ),
    .S0(_01546_),
    .S1(_01550_),
    .Z(_01873_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05385_ (.A1(_01554_),
    .A2(_01873_),
    .ZN(_01874_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05386_ (.I0(\u_cpu.rf_ram.memory[0][3] ),
    .I1(\u_cpu.rf_ram.memory[1][3] ),
    .I2(\u_cpu.rf_ram.memory[2][3] ),
    .I3(\u_cpu.rf_ram.memory[3][3] ),
    .S0(_01556_),
    .S1(_01557_),
    .Z(_01875_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05387_ (.A1(_01562_),
    .A2(_01875_),
    .B(_01565_),
    .ZN(_01876_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _05388_ (.A1(_01870_),
    .A2(_01872_),
    .B1(_01874_),
    .B2(_01876_),
    .C(_01568_),
    .ZN(_01877_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05389_ (.I0(\u_cpu.rf_ram.memory[20][3] ),
    .I1(\u_cpu.rf_ram.memory[21][3] ),
    .I2(\u_cpu.rf_ram.memory[22][3] ),
    .I3(\u_cpu.rf_ram.memory[23][3] ),
    .S0(_01572_),
    .S1(_01574_),
    .Z(_01878_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05390_ (.A1(_01570_),
    .A2(_01878_),
    .ZN(_01879_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05391_ (.I0(\u_cpu.rf_ram.memory[16][3] ),
    .I1(\u_cpu.rf_ram.memory[17][3] ),
    .I2(\u_cpu.rf_ram.memory[18][3] ),
    .I3(\u_cpu.rf_ram.memory[19][3] ),
    .S0(_01578_),
    .S1(_01580_),
    .Z(_01880_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05392_ (.A1(_01562_),
    .A2(_01880_),
    .B(_01582_),
    .ZN(_01881_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05393_ (.I0(\u_cpu.rf_ram.memory[28][3] ),
    .I1(\u_cpu.rf_ram.memory[29][3] ),
    .I2(\u_cpu.rf_ram.memory[30][3] ),
    .I3(\u_cpu.rf_ram.memory[31][3] ),
    .S0(_01572_),
    .S1(_01574_),
    .Z(_01882_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05394_ (.A1(_01570_),
    .A2(_01882_),
    .ZN(_01883_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05395_ (.I0(\u_cpu.rf_ram.memory[24][3] ),
    .I1(\u_cpu.rf_ram.memory[25][3] ),
    .I2(\u_cpu.rf_ram.memory[26][3] ),
    .I3(\u_cpu.rf_ram.memory[27][3] ),
    .S0(_01578_),
    .S1(_01580_),
    .Z(_01884_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05396_ (.A1(_01542_),
    .A2(_01884_),
    .B(_01418_),
    .ZN(_01885_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _05397_ (.A1(_01879_),
    .A2(_01881_),
    .B1(_01883_),
    .B2(_01885_),
    .C(_01426_),
    .ZN(_01886_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05398_ (.I0(\u_cpu.rf_ram.memory[52][3] ),
    .I1(\u_cpu.rf_ram.memory[53][3] ),
    .I2(\u_cpu.rf_ram.memory[54][3] ),
    .I3(\u_cpu.rf_ram.memory[55][3] ),
    .S0(_01590_),
    .S1(_01591_),
    .Z(_01887_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05399_ (.A1(_01589_),
    .A2(_01887_),
    .ZN(_01888_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05400_ (.I0(\u_cpu.rf_ram.memory[48][3] ),
    .I1(\u_cpu.rf_ram.memory[49][3] ),
    .I2(\u_cpu.rf_ram.memory[50][3] ),
    .I3(\u_cpu.rf_ram.memory[51][3] ),
    .S0(_01544_),
    .S1(_01548_),
    .Z(_01889_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05401_ (.A1(_01594_),
    .A2(_01889_),
    .B(_01564_),
    .ZN(_01890_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05402_ (.I0(\u_cpu.rf_ram.memory[60][3] ),
    .I1(\u_cpu.rf_ram.memory[61][3] ),
    .I2(\u_cpu.rf_ram.memory[62][3] ),
    .I3(\u_cpu.rf_ram.memory[63][3] ),
    .S0(_01598_),
    .S1(_01573_),
    .Z(_01891_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05403_ (.A1(_01597_),
    .A2(_01891_),
    .ZN(_01892_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05404_ (.I0(\u_cpu.rf_ram.memory[56][3] ),
    .I1(\u_cpu.rf_ram.memory[57][3] ),
    .I2(\u_cpu.rf_ram.memory[58][3] ),
    .I3(\u_cpu.rf_ram.memory[59][3] ),
    .S0(_01602_),
    .S1(_01579_),
    .Z(_01893_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05405_ (.A1(_01601_),
    .A2(_01893_),
    .B(_01605_),
    .ZN(_01894_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _05406_ (.A1(_01888_),
    .A2(_01890_),
    .B1(_01892_),
    .B2(_01894_),
    .C(_01607_),
    .ZN(_01895_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05407_ (.I0(\u_cpu.rf_ram.memory[40][3] ),
    .I1(\u_cpu.rf_ram.memory[41][3] ),
    .I2(\u_cpu.rf_ram.memory[42][3] ),
    .I3(\u_cpu.rf_ram.memory[43][3] ),
    .S0(_01545_),
    .S1(_01611_),
    .Z(_01896_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05408_ (.A1(_01609_),
    .A2(_01896_),
    .ZN(_01897_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05409_ (.I0(\u_cpu.rf_ram.memory[44][3] ),
    .I1(\u_cpu.rf_ram.memory[45][3] ),
    .I2(\u_cpu.rf_ram.memory[46][3] ),
    .I3(\u_cpu.rf_ram.memory[47][3] ),
    .S0(_01615_),
    .S1(_01616_),
    .Z(_01898_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05410_ (.A1(_01614_),
    .A2(_01898_),
    .B(_01605_),
    .ZN(_01899_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05411_ (.I0(\u_cpu.rf_ram.memory[36][3] ),
    .I1(\u_cpu.rf_ram.memory[37][3] ),
    .I2(\u_cpu.rf_ram.memory[38][3] ),
    .I3(\u_cpu.rf_ram.memory[39][3] ),
    .S0(_01619_),
    .S1(_01620_),
    .Z(_01900_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05412_ (.A1(_01589_),
    .A2(_01900_),
    .ZN(_01901_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05413_ (.I0(\u_cpu.rf_ram.memory[32][3] ),
    .I1(\u_cpu.rf_ram.memory[33][3] ),
    .I2(\u_cpu.rf_ram.memory[34][3] ),
    .I3(\u_cpu.rf_ram.memory[35][3] ),
    .S0(_01623_),
    .S1(_01624_),
    .Z(_01902_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05414_ (.A1(_01541_),
    .A2(_01902_),
    .B(_01626_),
    .ZN(_01903_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _05415_ (.A1(_01897_),
    .A2(_01899_),
    .B1(_01901_),
    .B2(_01903_),
    .C(_01628_),
    .ZN(_01904_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _05416_ (.A1(_01422_),
    .A2(_01895_),
    .A3(_01904_),
    .Z(_01905_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _05417_ (.A1(_01539_),
    .A2(_01877_),
    .A3(_01886_),
    .B(_01905_),
    .ZN(_01906_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05418_ (.I0(\u_cpu.rf_ram.memory[108][3] ),
    .I1(\u_cpu.rf_ram.memory[109][3] ),
    .I2(\u_cpu.rf_ram.memory[110][3] ),
    .I3(\u_cpu.rf_ram.memory[111][3] ),
    .S0(_01598_),
    .S1(_01573_),
    .Z(_01907_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05419_ (.A1(_01597_),
    .A2(_01907_),
    .ZN(_01908_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05420_ (.I0(\u_cpu.rf_ram.memory[104][3] ),
    .I1(\u_cpu.rf_ram.memory[105][3] ),
    .I2(\u_cpu.rf_ram.memory[106][3] ),
    .I3(\u_cpu.rf_ram.memory[107][3] ),
    .S0(_01615_),
    .S1(_01616_),
    .Z(_01909_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05421_ (.A1(_01594_),
    .A2(_01909_),
    .B(_01416_),
    .ZN(_01910_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05422_ (.I0(\u_cpu.rf_ram.memory[100][3] ),
    .I1(\u_cpu.rf_ram.memory[101][3] ),
    .I2(\u_cpu.rf_ram.memory[102][3] ),
    .I3(\u_cpu.rf_ram.memory[103][3] ),
    .S0(_01577_),
    .S1(_01549_),
    .Z(_01911_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05423_ (.A1(_01636_),
    .A2(_01911_),
    .ZN(_01912_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05424_ (.I0(\u_cpu.rf_ram.memory[96][3] ),
    .I1(\u_cpu.rf_ram.memory[97][3] ),
    .I2(\u_cpu.rf_ram.memory[98][3] ),
    .I3(\u_cpu.rf_ram.memory[99][3] ),
    .S0(_01602_),
    .S1(_01579_),
    .Z(_01913_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05425_ (.A1(_01601_),
    .A2(_01913_),
    .B(_01626_),
    .ZN(_01914_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _05426_ (.A1(_01908_),
    .A2(_01910_),
    .B1(_01912_),
    .B2(_01914_),
    .C(_01628_),
    .ZN(_01915_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05427_ (.I0(\u_cpu.rf_ram.memory[124][3] ),
    .I1(\u_cpu.rf_ram.memory[125][3] ),
    .I2(\u_cpu.rf_ram.memory[126][3] ),
    .I3(\u_cpu.rf_ram.memory[127][3] ),
    .S0(_01545_),
    .S1(_01642_),
    .Z(_01916_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05428_ (.A1(_01398_),
    .A2(_01916_),
    .ZN(_01917_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05429_ (.I0(\u_cpu.rf_ram.memory[120][3] ),
    .I1(\u_cpu.rf_ram.memory[121][3] ),
    .I2(\u_cpu.rf_ram.memory[122][3] ),
    .I3(\u_cpu.rf_ram.memory[123][3] ),
    .S0(_01646_),
    .S1(_01603_),
    .Z(_01918_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05430_ (.A1(_01645_),
    .A2(_01918_),
    .B(_01648_),
    .ZN(_01919_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05431_ (.I0(\u_cpu.rf_ram.memory[112][3] ),
    .I1(\u_cpu.rf_ram.memory[113][3] ),
    .I2(\u_cpu.rf_ram.memory[114][3] ),
    .I3(\u_cpu.rf_ram.memory[115][3] ),
    .S0(_01619_),
    .S1(_01620_),
    .Z(_01920_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05432_ (.A1(_01541_),
    .A2(_01920_),
    .ZN(_01921_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05433_ (.I0(\u_cpu.rf_ram.memory[116][3] ),
    .I1(\u_cpu.rf_ram.memory[117][3] ),
    .I2(\u_cpu.rf_ram.memory[118][3] ),
    .I3(\u_cpu.rf_ram.memory[119][3] ),
    .S0(_01623_),
    .S1(_01624_),
    .Z(_01922_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05434_ (.A1(_01614_),
    .A2(_01922_),
    .B(_01654_),
    .ZN(_01923_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _05435_ (.A1(_01917_),
    .A2(_01919_),
    .B1(_01921_),
    .B2(_01923_),
    .C(_01607_),
    .ZN(_01924_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _05436_ (.A1(_01422_),
    .A2(_01915_),
    .A3(_01924_),
    .ZN(_01925_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05437_ (.I0(\u_cpu.rf_ram.memory[92][3] ),
    .I1(\u_cpu.rf_ram.memory[93][3] ),
    .I2(\u_cpu.rf_ram.memory[94][3] ),
    .I3(\u_cpu.rf_ram.memory[95][3] ),
    .S0(_01610_),
    .S1(_01611_),
    .Z(_01926_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05438_ (.A1(_01398_),
    .A2(_01926_),
    .ZN(_01927_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05439_ (.I0(\u_cpu.rf_ram.memory[88][3] ),
    .I1(\u_cpu.rf_ram.memory[89][3] ),
    .I2(\u_cpu.rf_ram.memory[90][3] ),
    .I3(\u_cpu.rf_ram.memory[91][3] ),
    .S0(_01646_),
    .S1(_01603_),
    .Z(_01928_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05440_ (.A1(_01645_),
    .A2(_01928_),
    .B(_01648_),
    .ZN(_01929_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05441_ (.I0(\u_cpu.rf_ram.memory[80][3] ),
    .I1(\u_cpu.rf_ram.memory[81][3] ),
    .I2(\u_cpu.rf_ram.memory[82][3] ),
    .I3(\u_cpu.rf_ram.memory[83][3] ),
    .S0(_01590_),
    .S1(_01642_),
    .Z(_01930_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05442_ (.A1(_01609_),
    .A2(_01930_),
    .ZN(_01931_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05443_ (.I0(\u_cpu.rf_ram.memory[84][3] ),
    .I1(\u_cpu.rf_ram.memory[85][3] ),
    .I2(\u_cpu.rf_ram.memory[86][3] ),
    .I3(\u_cpu.rf_ram.memory[87][3] ),
    .S0(_01555_),
    .S1(_01652_),
    .Z(_01932_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05444_ (.A1(_01553_),
    .A2(_01932_),
    .B(_01654_),
    .ZN(_01933_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _05445_ (.A1(_01927_),
    .A2(_01929_),
    .B1(_01931_),
    .B2(_01933_),
    .C(_01426_),
    .ZN(_01934_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05446_ (.I0(\u_cpu.rf_ram.memory[64][3] ),
    .I1(\u_cpu.rf_ram.memory[65][3] ),
    .I2(\u_cpu.rf_ram.memory[66][3] ),
    .I3(\u_cpu.rf_ram.memory[67][3] ),
    .S0(_01571_),
    .S1(_01668_),
    .Z(_01935_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05447_ (.A1(_01667_),
    .A2(_01935_),
    .ZN(_01936_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05448_ (.I0(\u_cpu.rf_ram.memory[68][3] ),
    .I1(\u_cpu.rf_ram.memory[69][3] ),
    .I2(\u_cpu.rf_ram.memory[70][3] ),
    .I3(\u_cpu.rf_ram.memory[71][3] ),
    .S0(_01555_),
    .S1(_01652_),
    .Z(_01937_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05449_ (.A1(_01553_),
    .A2(_01937_),
    .B(_01565_),
    .ZN(_01938_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05450_ (.I0(\u_cpu.rf_ram.memory[72][3] ),
    .I1(\u_cpu.rf_ram.memory[73][3] ),
    .I2(\u_cpu.rf_ram.memory[74][3] ),
    .I3(\u_cpu.rf_ram.memory[75][3] ),
    .S0(_01610_),
    .S1(_01668_),
    .Z(_01939_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05451_ (.A1(_01667_),
    .A2(_01939_),
    .ZN(_01940_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05452_ (.I0(\u_cpu.rf_ram.memory[76][3] ),
    .I1(\u_cpu.rf_ram.memory[77][3] ),
    .I2(\u_cpu.rf_ram.memory[78][3] ),
    .I3(\u_cpu.rf_ram.memory[79][3] ),
    .S0(_01577_),
    .S1(_01549_),
    .Z(_01941_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05453_ (.A1(_01636_),
    .A2(_01941_),
    .B(_01417_),
    .ZN(_01942_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _05454_ (.A1(_01936_),
    .A2(_01938_),
    .B1(_01940_),
    .B2(_01942_),
    .C(_01568_),
    .ZN(_01943_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _05455_ (.A1(_01539_),
    .A2(_01934_),
    .A3(_01943_),
    .ZN(_01944_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05456_ (.A1(_01925_),
    .A2(_01944_),
    .B(_01402_),
    .ZN(_01945_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05457_ (.I0(\u_cpu.rf_ram.memory[136][3] ),
    .I1(\u_cpu.rf_ram.memory[137][3] ),
    .I2(\u_cpu.rf_ram.memory[138][3] ),
    .I3(\u_cpu.rf_ram.memory[139][3] ),
    .S0(_01680_),
    .S1(_01681_),
    .Z(_01946_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05458_ (.A1(_01399_),
    .A2(_01946_),
    .ZN(_01947_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05459_ (.I0(\u_cpu.rf_ram.memory[140][3] ),
    .I1(\u_cpu.rf_ram.memory[141][3] ),
    .I2(\u_cpu.rf_ram.memory[142][3] ),
    .I3(\u_cpu.rf_ram.memory[143][3] ),
    .S0(_01680_),
    .S1(_01681_),
    .Z(_01948_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05460_ (.A1(_01684_),
    .A2(_01948_),
    .B(_01582_),
    .ZN(_01949_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05461_ (.I0(\u_cpu.rf_ram.memory[128][3] ),
    .I1(\u_cpu.rf_ram.memory[129][3] ),
    .I2(\u_cpu.rf_ram.memory[130][3] ),
    .I3(\u_cpu.rf_ram.memory[131][3] ),
    .S0(_01687_),
    .S1(_01688_),
    .Z(_01950_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05462_ (.A1(_01399_),
    .A2(_01950_),
    .ZN(_01951_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05463_ (.I0(\u_cpu.rf_ram.memory[132][3] ),
    .I1(\u_cpu.rf_ram.memory[133][3] ),
    .I2(\u_cpu.rf_ram.memory[134][3] ),
    .I3(\u_cpu.rf_ram.memory[135][3] ),
    .S0(_01687_),
    .S1(_01688_),
    .Z(_01952_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05464_ (.A1(_01684_),
    .A2(_01952_),
    .B(_01418_),
    .ZN(_01953_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _05465_ (.A1(_01947_),
    .A2(_01949_),
    .B1(_01951_),
    .B2(_01953_),
    .C(_01404_),
    .ZN(_01954_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05466_ (.A1(_01945_),
    .A2(_01954_),
    .ZN(_01955_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05467_ (.A1(_01406_),
    .A2(_01906_),
    .B(_01955_),
    .ZN(_00003_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05468_ (.I0(\u_cpu.rf_ram.memory[8][4] ),
    .I1(\u_cpu.rf_ram.memory[9][4] ),
    .I2(\u_cpu.rf_ram.memory[10][4] ),
    .I3(\u_cpu.rf_ram.memory[11][4] ),
    .S0(_01546_),
    .S1(_01550_),
    .Z(_01956_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05469_ (.A1(_01542_),
    .A2(_01956_),
    .ZN(_01957_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05470_ (.I0(\u_cpu.rf_ram.memory[12][4] ),
    .I1(\u_cpu.rf_ram.memory[13][4] ),
    .I2(\u_cpu.rf_ram.memory[14][4] ),
    .I3(\u_cpu.rf_ram.memory[15][4] ),
    .S0(_01556_),
    .S1(_01557_),
    .Z(_01958_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05471_ (.A1(_01554_),
    .A2(_01958_),
    .B(_01417_),
    .ZN(_01959_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05472_ (.I0(\u_cpu.rf_ram.memory[4][4] ),
    .I1(\u_cpu.rf_ram.memory[5][4] ),
    .I2(\u_cpu.rf_ram.memory[6][4] ),
    .I3(\u_cpu.rf_ram.memory[7][4] ),
    .S0(_01546_),
    .S1(_01550_),
    .Z(_01960_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05473_ (.A1(_01554_),
    .A2(_01960_),
    .ZN(_01961_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05474_ (.I0(\u_cpu.rf_ram.memory[0][4] ),
    .I1(\u_cpu.rf_ram.memory[1][4] ),
    .I2(\u_cpu.rf_ram.memory[2][4] ),
    .I3(\u_cpu.rf_ram.memory[3][4] ),
    .S0(_01556_),
    .S1(_01557_),
    .Z(_01962_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05475_ (.A1(_01562_),
    .A2(_01962_),
    .B(_01565_),
    .ZN(_01963_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _05476_ (.A1(_01957_),
    .A2(_01959_),
    .B1(_01961_),
    .B2(_01963_),
    .C(_01568_),
    .ZN(_01964_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05477_ (.I0(\u_cpu.rf_ram.memory[20][4] ),
    .I1(\u_cpu.rf_ram.memory[21][4] ),
    .I2(\u_cpu.rf_ram.memory[22][4] ),
    .I3(\u_cpu.rf_ram.memory[23][4] ),
    .S0(_01572_),
    .S1(_01574_),
    .Z(_01965_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05478_ (.A1(_01570_),
    .A2(_01965_),
    .ZN(_01966_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05479_ (.I0(\u_cpu.rf_ram.memory[16][4] ),
    .I1(\u_cpu.rf_ram.memory[17][4] ),
    .I2(\u_cpu.rf_ram.memory[18][4] ),
    .I3(\u_cpu.rf_ram.memory[19][4] ),
    .S0(_01578_),
    .S1(_01580_),
    .Z(_01967_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05480_ (.A1(_01562_),
    .A2(_01967_),
    .B(_01582_),
    .ZN(_01968_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05481_ (.I0(\u_cpu.rf_ram.memory[28][4] ),
    .I1(\u_cpu.rf_ram.memory[29][4] ),
    .I2(\u_cpu.rf_ram.memory[30][4] ),
    .I3(\u_cpu.rf_ram.memory[31][4] ),
    .S0(_01572_),
    .S1(_01574_),
    .Z(_01969_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05482_ (.A1(_01570_),
    .A2(_01969_),
    .ZN(_01970_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05483_ (.I0(\u_cpu.rf_ram.memory[24][4] ),
    .I1(\u_cpu.rf_ram.memory[25][4] ),
    .I2(\u_cpu.rf_ram.memory[26][4] ),
    .I3(\u_cpu.rf_ram.memory[27][4] ),
    .S0(_01578_),
    .S1(_01580_),
    .Z(_01971_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05484_ (.A1(_01542_),
    .A2(_01971_),
    .B(_01418_),
    .ZN(_01972_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _05485_ (.A1(_01966_),
    .A2(_01968_),
    .B1(_01970_),
    .B2(_01972_),
    .C(_01426_),
    .ZN(_01973_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05486_ (.I0(\u_cpu.rf_ram.memory[52][4] ),
    .I1(\u_cpu.rf_ram.memory[53][4] ),
    .I2(\u_cpu.rf_ram.memory[54][4] ),
    .I3(\u_cpu.rf_ram.memory[55][4] ),
    .S0(_01590_),
    .S1(_01591_),
    .Z(_01974_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05487_ (.A1(_01589_),
    .A2(_01974_),
    .ZN(_01975_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05488_ (.I0(\u_cpu.rf_ram.memory[48][4] ),
    .I1(\u_cpu.rf_ram.memory[49][4] ),
    .I2(\u_cpu.rf_ram.memory[50][4] ),
    .I3(\u_cpu.rf_ram.memory[51][4] ),
    .S0(_01544_),
    .S1(_01548_),
    .Z(_01976_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05489_ (.A1(_01594_),
    .A2(_01976_),
    .B(_01564_),
    .ZN(_01977_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05490_ (.I0(\u_cpu.rf_ram.memory[60][4] ),
    .I1(\u_cpu.rf_ram.memory[61][4] ),
    .I2(\u_cpu.rf_ram.memory[62][4] ),
    .I3(\u_cpu.rf_ram.memory[63][4] ),
    .S0(_01598_),
    .S1(_01573_),
    .Z(_01978_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05491_ (.A1(_01597_),
    .A2(_01978_),
    .ZN(_01979_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05492_ (.I0(\u_cpu.rf_ram.memory[56][4] ),
    .I1(\u_cpu.rf_ram.memory[57][4] ),
    .I2(\u_cpu.rf_ram.memory[58][4] ),
    .I3(\u_cpu.rf_ram.memory[59][4] ),
    .S0(_01602_),
    .S1(_01579_),
    .Z(_01980_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05493_ (.A1(_01601_),
    .A2(_01980_),
    .B(_01605_),
    .ZN(_01981_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _05494_ (.A1(_01975_),
    .A2(_01977_),
    .B1(_01979_),
    .B2(_01981_),
    .C(_01607_),
    .ZN(_01982_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05495_ (.I0(\u_cpu.rf_ram.memory[40][4] ),
    .I1(\u_cpu.rf_ram.memory[41][4] ),
    .I2(\u_cpu.rf_ram.memory[42][4] ),
    .I3(\u_cpu.rf_ram.memory[43][4] ),
    .S0(_01545_),
    .S1(_01642_),
    .Z(_01983_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05496_ (.A1(_01609_),
    .A2(_01983_),
    .ZN(_01984_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05497_ (.I0(\u_cpu.rf_ram.memory[44][4] ),
    .I1(\u_cpu.rf_ram.memory[45][4] ),
    .I2(\u_cpu.rf_ram.memory[46][4] ),
    .I3(\u_cpu.rf_ram.memory[47][4] ),
    .S0(_01615_),
    .S1(_01616_),
    .Z(_01985_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05498_ (.A1(_01397_),
    .A2(_01985_),
    .B(_01605_),
    .ZN(_01986_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05499_ (.I0(\u_cpu.rf_ram.memory[36][4] ),
    .I1(\u_cpu.rf_ram.memory[37][4] ),
    .I2(\u_cpu.rf_ram.memory[38][4] ),
    .I3(\u_cpu.rf_ram.memory[39][4] ),
    .S0(_01619_),
    .S1(_01620_),
    .Z(_01987_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05500_ (.A1(_01589_),
    .A2(_01987_),
    .ZN(_01988_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05501_ (.I0(\u_cpu.rf_ram.memory[32][4] ),
    .I1(\u_cpu.rf_ram.memory[33][4] ),
    .I2(\u_cpu.rf_ram.memory[34][4] ),
    .I3(\u_cpu.rf_ram.memory[35][4] ),
    .S0(_01623_),
    .S1(_01624_),
    .Z(_01989_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05502_ (.A1(_01541_),
    .A2(_01989_),
    .B(_01626_),
    .ZN(_01990_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _05503_ (.A1(_01984_),
    .A2(_01986_),
    .B1(_01988_),
    .B2(_01990_),
    .C(_01628_),
    .ZN(_01991_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _05504_ (.A1(_01422_),
    .A2(_01982_),
    .A3(_01991_),
    .Z(_01992_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _05505_ (.A1(_01539_),
    .A2(_01964_),
    .A3(_01973_),
    .B(_01992_),
    .ZN(_01993_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05506_ (.I0(\u_cpu.rf_ram.memory[108][4] ),
    .I1(\u_cpu.rf_ram.memory[109][4] ),
    .I2(\u_cpu.rf_ram.memory[110][4] ),
    .I3(\u_cpu.rf_ram.memory[111][4] ),
    .S0(_01598_),
    .S1(_01573_),
    .Z(_01994_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05507_ (.A1(_01597_),
    .A2(_01994_),
    .ZN(_01995_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05508_ (.I0(\u_cpu.rf_ram.memory[104][4] ),
    .I1(\u_cpu.rf_ram.memory[105][4] ),
    .I2(\u_cpu.rf_ram.memory[106][4] ),
    .I3(\u_cpu.rf_ram.memory[107][4] ),
    .S0(_01615_),
    .S1(_01616_),
    .Z(_01996_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05509_ (.A1(_01594_),
    .A2(_01996_),
    .B(_01416_),
    .ZN(_01997_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05510_ (.I0(\u_cpu.rf_ram.memory[100][4] ),
    .I1(\u_cpu.rf_ram.memory[101][4] ),
    .I2(\u_cpu.rf_ram.memory[102][4] ),
    .I3(\u_cpu.rf_ram.memory[103][4] ),
    .S0(_01577_),
    .S1(_01549_),
    .Z(_01998_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05511_ (.A1(_01636_),
    .A2(_01998_),
    .ZN(_01999_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05512_ (.I0(\u_cpu.rf_ram.memory[96][4] ),
    .I1(\u_cpu.rf_ram.memory[97][4] ),
    .I2(\u_cpu.rf_ram.memory[98][4] ),
    .I3(\u_cpu.rf_ram.memory[99][4] ),
    .S0(_01602_),
    .S1(_01579_),
    .Z(_02000_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05513_ (.A1(_01601_),
    .A2(_02000_),
    .B(_01626_),
    .ZN(_02001_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _05514_ (.A1(_01995_),
    .A2(_01997_),
    .B1(_01999_),
    .B2(_02001_),
    .C(_01628_),
    .ZN(_02002_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05515_ (.I0(\u_cpu.rf_ram.memory[124][4] ),
    .I1(\u_cpu.rf_ram.memory[125][4] ),
    .I2(\u_cpu.rf_ram.memory[126][4] ),
    .I3(\u_cpu.rf_ram.memory[127][4] ),
    .S0(_01545_),
    .S1(_01642_),
    .Z(_02003_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05516_ (.A1(_01398_),
    .A2(_02003_),
    .ZN(_02004_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05517_ (.I0(\u_cpu.rf_ram.memory[120][4] ),
    .I1(\u_cpu.rf_ram.memory[121][4] ),
    .I2(\u_cpu.rf_ram.memory[122][4] ),
    .I3(\u_cpu.rf_ram.memory[123][4] ),
    .S0(_01646_),
    .S1(_01603_),
    .Z(_02005_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05518_ (.A1(_01645_),
    .A2(_02005_),
    .B(_01648_),
    .ZN(_02006_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05519_ (.I0(\u_cpu.rf_ram.memory[112][4] ),
    .I1(\u_cpu.rf_ram.memory[113][4] ),
    .I2(\u_cpu.rf_ram.memory[114][4] ),
    .I3(\u_cpu.rf_ram.memory[115][4] ),
    .S0(_01619_),
    .S1(_01620_),
    .Z(_02007_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05520_ (.A1(_01541_),
    .A2(_02007_),
    .ZN(_02008_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05521_ (.I0(\u_cpu.rf_ram.memory[116][4] ),
    .I1(\u_cpu.rf_ram.memory[117][4] ),
    .I2(\u_cpu.rf_ram.memory[118][4] ),
    .I3(\u_cpu.rf_ram.memory[119][4] ),
    .S0(_01623_),
    .S1(_01624_),
    .Z(_02009_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05522_ (.A1(_01614_),
    .A2(_02009_),
    .B(_01654_),
    .ZN(_02010_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _05523_ (.A1(_02004_),
    .A2(_02006_),
    .B1(_02008_),
    .B2(_02010_),
    .C(_01607_),
    .ZN(_02011_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _05524_ (.A1(_01422_),
    .A2(_02002_),
    .A3(_02011_),
    .ZN(_02012_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05525_ (.I0(\u_cpu.rf_ram.memory[92][4] ),
    .I1(\u_cpu.rf_ram.memory[93][4] ),
    .I2(\u_cpu.rf_ram.memory[94][4] ),
    .I3(\u_cpu.rf_ram.memory[95][4] ),
    .S0(_01610_),
    .S1(_01611_),
    .Z(_02013_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05526_ (.A1(_01398_),
    .A2(_02013_),
    .ZN(_02014_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05527_ (.I0(\u_cpu.rf_ram.memory[88][4] ),
    .I1(\u_cpu.rf_ram.memory[89][4] ),
    .I2(\u_cpu.rf_ram.memory[90][4] ),
    .I3(\u_cpu.rf_ram.memory[91][4] ),
    .S0(_01646_),
    .S1(_01603_),
    .Z(_02015_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05528_ (.A1(_01645_),
    .A2(_02015_),
    .B(_01648_),
    .ZN(_02016_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05529_ (.I0(\u_cpu.rf_ram.memory[80][4] ),
    .I1(\u_cpu.rf_ram.memory[81][4] ),
    .I2(\u_cpu.rf_ram.memory[82][4] ),
    .I3(\u_cpu.rf_ram.memory[83][4] ),
    .S0(_01590_),
    .S1(_01591_),
    .Z(_02017_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05530_ (.A1(_01609_),
    .A2(_02017_),
    .ZN(_02018_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05531_ (.I0(\u_cpu.rf_ram.memory[84][4] ),
    .I1(\u_cpu.rf_ram.memory[85][4] ),
    .I2(\u_cpu.rf_ram.memory[86][4] ),
    .I3(\u_cpu.rf_ram.memory[87][4] ),
    .S0(_01555_),
    .S1(_01652_),
    .Z(_02019_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05532_ (.A1(_01614_),
    .A2(_02019_),
    .B(_01654_),
    .ZN(_02020_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _05533_ (.A1(_02014_),
    .A2(_02016_),
    .B1(_02018_),
    .B2(_02020_),
    .C(_01426_),
    .ZN(_02021_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05534_ (.I0(\u_cpu.rf_ram.memory[64][4] ),
    .I1(\u_cpu.rf_ram.memory[65][4] ),
    .I2(\u_cpu.rf_ram.memory[66][4] ),
    .I3(\u_cpu.rf_ram.memory[67][4] ),
    .S0(_01571_),
    .S1(_01668_),
    .Z(_02022_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05535_ (.A1(_01667_),
    .A2(_02022_),
    .ZN(_02023_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05536_ (.I0(\u_cpu.rf_ram.memory[68][4] ),
    .I1(\u_cpu.rf_ram.memory[69][4] ),
    .I2(\u_cpu.rf_ram.memory[70][4] ),
    .I3(\u_cpu.rf_ram.memory[71][4] ),
    .S0(_01555_),
    .S1(_01652_),
    .Z(_02024_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05537_ (.A1(_01553_),
    .A2(_02024_),
    .B(_01565_),
    .ZN(_02025_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05538_ (.I0(\u_cpu.rf_ram.memory[72][4] ),
    .I1(\u_cpu.rf_ram.memory[73][4] ),
    .I2(\u_cpu.rf_ram.memory[74][4] ),
    .I3(\u_cpu.rf_ram.memory[75][4] ),
    .S0(_01610_),
    .S1(_01611_),
    .Z(_02026_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05539_ (.A1(_01667_),
    .A2(_02026_),
    .ZN(_02027_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05540_ (.I0(\u_cpu.rf_ram.memory[76][4] ),
    .I1(\u_cpu.rf_ram.memory[77][4] ),
    .I2(\u_cpu.rf_ram.memory[78][4] ),
    .I3(\u_cpu.rf_ram.memory[79][4] ),
    .S0(_01577_),
    .S1(_01549_),
    .Z(_02028_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05541_ (.A1(_01636_),
    .A2(_02028_),
    .B(_01417_),
    .ZN(_02029_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _05542_ (.A1(_02023_),
    .A2(_02025_),
    .B1(_02027_),
    .B2(_02029_),
    .C(_01568_),
    .ZN(_02030_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _05543_ (.A1(_01539_),
    .A2(_02021_),
    .A3(_02030_),
    .ZN(_02031_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05544_ (.A1(_02012_),
    .A2(_02031_),
    .B(_01402_),
    .ZN(_02032_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05545_ (.I0(\u_cpu.rf_ram.memory[136][4] ),
    .I1(\u_cpu.rf_ram.memory[137][4] ),
    .I2(\u_cpu.rf_ram.memory[138][4] ),
    .I3(\u_cpu.rf_ram.memory[139][4] ),
    .S0(_01680_),
    .S1(_01681_),
    .Z(_02033_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05546_ (.A1(_01399_),
    .A2(_02033_),
    .ZN(_02034_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05547_ (.I0(\u_cpu.rf_ram.memory[140][4] ),
    .I1(\u_cpu.rf_ram.memory[141][4] ),
    .I2(\u_cpu.rf_ram.memory[142][4] ),
    .I3(\u_cpu.rf_ram.memory[143][4] ),
    .S0(_01680_),
    .S1(_01681_),
    .Z(_02035_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05548_ (.A1(_01684_),
    .A2(_02035_),
    .B(_01582_),
    .ZN(_02036_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05549_ (.I0(\u_cpu.rf_ram.memory[128][4] ),
    .I1(\u_cpu.rf_ram.memory[129][4] ),
    .I2(\u_cpu.rf_ram.memory[130][4] ),
    .I3(\u_cpu.rf_ram.memory[131][4] ),
    .S0(_01687_),
    .S1(_01688_),
    .Z(_02037_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05550_ (.A1(_01399_),
    .A2(_02037_),
    .ZN(_02038_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05551_ (.I0(\u_cpu.rf_ram.memory[132][4] ),
    .I1(\u_cpu.rf_ram.memory[133][4] ),
    .I2(\u_cpu.rf_ram.memory[134][4] ),
    .I3(\u_cpu.rf_ram.memory[135][4] ),
    .S0(_01687_),
    .S1(_01688_),
    .Z(_02039_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05552_ (.A1(_01684_),
    .A2(_02039_),
    .B(_01418_),
    .ZN(_02040_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _05553_ (.A1(_02034_),
    .A2(_02036_),
    .B1(_02038_),
    .B2(_02040_),
    .C(_01404_),
    .ZN(_02041_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05554_ (.A1(_02032_),
    .A2(_02041_),
    .ZN(_02042_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05555_ (.A1(_01406_),
    .A2(_01993_),
    .B(_02042_),
    .ZN(_00004_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05556_ (.I0(\u_cpu.rf_ram.memory[8][5] ),
    .I1(\u_cpu.rf_ram.memory[9][5] ),
    .I2(\u_cpu.rf_ram.memory[10][5] ),
    .I3(\u_cpu.rf_ram.memory[11][5] ),
    .S0(_01546_),
    .S1(_01550_),
    .Z(_02043_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05557_ (.A1(_01542_),
    .A2(_02043_),
    .ZN(_02044_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05558_ (.I0(\u_cpu.rf_ram.memory[12][5] ),
    .I1(\u_cpu.rf_ram.memory[13][5] ),
    .I2(\u_cpu.rf_ram.memory[14][5] ),
    .I3(\u_cpu.rf_ram.memory[15][5] ),
    .S0(_01556_),
    .S1(_01557_),
    .Z(_02045_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05559_ (.A1(_01554_),
    .A2(_02045_),
    .B(_01417_),
    .ZN(_02046_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05560_ (.I0(\u_cpu.rf_ram.memory[4][5] ),
    .I1(\u_cpu.rf_ram.memory[5][5] ),
    .I2(\u_cpu.rf_ram.memory[6][5] ),
    .I3(\u_cpu.rf_ram.memory[7][5] ),
    .S0(_01546_),
    .S1(_01550_),
    .Z(_02047_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05561_ (.A1(_01554_),
    .A2(_02047_),
    .ZN(_02048_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05562_ (.I0(\u_cpu.rf_ram.memory[0][5] ),
    .I1(\u_cpu.rf_ram.memory[1][5] ),
    .I2(\u_cpu.rf_ram.memory[2][5] ),
    .I3(\u_cpu.rf_ram.memory[3][5] ),
    .S0(_01556_),
    .S1(_01557_),
    .Z(_02049_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05563_ (.A1(_01562_),
    .A2(_02049_),
    .B(_01565_),
    .ZN(_02050_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _05564_ (.A1(_02044_),
    .A2(_02046_),
    .B1(_02048_),
    .B2(_02050_),
    .C(_01568_),
    .ZN(_02051_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05565_ (.I0(\u_cpu.rf_ram.memory[20][5] ),
    .I1(\u_cpu.rf_ram.memory[21][5] ),
    .I2(\u_cpu.rf_ram.memory[22][5] ),
    .I3(\u_cpu.rf_ram.memory[23][5] ),
    .S0(_01572_),
    .S1(_01574_),
    .Z(_02052_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05566_ (.A1(_01570_),
    .A2(_02052_),
    .ZN(_02053_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05567_ (.I0(\u_cpu.rf_ram.memory[16][5] ),
    .I1(\u_cpu.rf_ram.memory[17][5] ),
    .I2(\u_cpu.rf_ram.memory[18][5] ),
    .I3(\u_cpu.rf_ram.memory[19][5] ),
    .S0(_01578_),
    .S1(_01580_),
    .Z(_02054_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05568_ (.A1(_01562_),
    .A2(_02054_),
    .B(_01582_),
    .ZN(_02055_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05569_ (.I0(\u_cpu.rf_ram.memory[28][5] ),
    .I1(\u_cpu.rf_ram.memory[29][5] ),
    .I2(\u_cpu.rf_ram.memory[30][5] ),
    .I3(\u_cpu.rf_ram.memory[31][5] ),
    .S0(_01572_),
    .S1(_01574_),
    .Z(_02056_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05570_ (.A1(_01570_),
    .A2(_02056_),
    .ZN(_02057_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05571_ (.I0(\u_cpu.rf_ram.memory[24][5] ),
    .I1(\u_cpu.rf_ram.memory[25][5] ),
    .I2(\u_cpu.rf_ram.memory[26][5] ),
    .I3(\u_cpu.rf_ram.memory[27][5] ),
    .S0(_01578_),
    .S1(_01580_),
    .Z(_02058_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05572_ (.A1(_01542_),
    .A2(_02058_),
    .B(_01418_),
    .ZN(_02059_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _05573_ (.A1(_02053_),
    .A2(_02055_),
    .B1(_02057_),
    .B2(_02059_),
    .C(_01426_),
    .ZN(_02060_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05574_ (.I0(\u_cpu.rf_ram.memory[52][5] ),
    .I1(\u_cpu.rf_ram.memory[53][5] ),
    .I2(\u_cpu.rf_ram.memory[54][5] ),
    .I3(\u_cpu.rf_ram.memory[55][5] ),
    .S0(_01590_),
    .S1(_01591_),
    .Z(_02061_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05575_ (.A1(_01589_),
    .A2(_02061_),
    .ZN(_02062_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05576_ (.I0(\u_cpu.rf_ram.memory[48][5] ),
    .I1(\u_cpu.rf_ram.memory[49][5] ),
    .I2(\u_cpu.rf_ram.memory[50][5] ),
    .I3(\u_cpu.rf_ram.memory[51][5] ),
    .S0(_01544_),
    .S1(_01548_),
    .Z(_02063_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05577_ (.A1(_01540_),
    .A2(_02063_),
    .B(_01564_),
    .ZN(_02064_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05578_ (.I0(\u_cpu.rf_ram.memory[60][5] ),
    .I1(\u_cpu.rf_ram.memory[61][5] ),
    .I2(\u_cpu.rf_ram.memory[62][5] ),
    .I3(\u_cpu.rf_ram.memory[63][5] ),
    .S0(_01598_),
    .S1(_01573_),
    .Z(_02065_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05579_ (.A1(_01636_),
    .A2(_02065_),
    .ZN(_02066_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05580_ (.I0(\u_cpu.rf_ram.memory[56][5] ),
    .I1(\u_cpu.rf_ram.memory[57][5] ),
    .I2(\u_cpu.rf_ram.memory[58][5] ),
    .I3(\u_cpu.rf_ram.memory[59][5] ),
    .S0(_01602_),
    .S1(_01579_),
    .Z(_02067_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05581_ (.A1(_01601_),
    .A2(_02067_),
    .B(_01605_),
    .ZN(_02068_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _05582_ (.A1(_02062_),
    .A2(_02064_),
    .B1(_02066_),
    .B2(_02068_),
    .C(_01607_),
    .ZN(_02069_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05583_ (.I0(\u_cpu.rf_ram.memory[40][5] ),
    .I1(\u_cpu.rf_ram.memory[41][5] ),
    .I2(\u_cpu.rf_ram.memory[42][5] ),
    .I3(\u_cpu.rf_ram.memory[43][5] ),
    .S0(_01545_),
    .S1(_01642_),
    .Z(_02070_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05584_ (.A1(_01609_),
    .A2(_02070_),
    .ZN(_02071_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05585_ (.I0(\u_cpu.rf_ram.memory[44][5] ),
    .I1(\u_cpu.rf_ram.memory[45][5] ),
    .I2(\u_cpu.rf_ram.memory[46][5] ),
    .I3(\u_cpu.rf_ram.memory[47][5] ),
    .S0(_01615_),
    .S1(_01616_),
    .Z(_02072_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05586_ (.A1(_01397_),
    .A2(_02072_),
    .B(_01605_),
    .ZN(_02073_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05587_ (.I0(\u_cpu.rf_ram.memory[36][5] ),
    .I1(\u_cpu.rf_ram.memory[37][5] ),
    .I2(\u_cpu.rf_ram.memory[38][5] ),
    .I3(\u_cpu.rf_ram.memory[39][5] ),
    .S0(_01619_),
    .S1(_01620_),
    .Z(_02074_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05588_ (.A1(_01597_),
    .A2(_02074_),
    .ZN(_02075_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05589_ (.I0(\u_cpu.rf_ram.memory[32][5] ),
    .I1(\u_cpu.rf_ram.memory[33][5] ),
    .I2(\u_cpu.rf_ram.memory[34][5] ),
    .I3(\u_cpu.rf_ram.memory[35][5] ),
    .S0(_01623_),
    .S1(_01624_),
    .Z(_02076_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05590_ (.A1(_01645_),
    .A2(_02076_),
    .B(_01626_),
    .ZN(_02077_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _05591_ (.A1(_02071_),
    .A2(_02073_),
    .B1(_02075_),
    .B2(_02077_),
    .C(_01628_),
    .ZN(_02078_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _05592_ (.A1(_01422_),
    .A2(_02069_),
    .A3(_02078_),
    .Z(_02079_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _05593_ (.A1(_01539_),
    .A2(_02051_),
    .A3(_02060_),
    .B(_02079_),
    .ZN(_02080_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05594_ (.I0(\u_cpu.rf_ram.memory[108][5] ),
    .I1(\u_cpu.rf_ram.memory[109][5] ),
    .I2(\u_cpu.rf_ram.memory[110][5] ),
    .I3(\u_cpu.rf_ram.memory[111][5] ),
    .S0(_01598_),
    .S1(_01573_),
    .Z(_02081_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05595_ (.A1(_01597_),
    .A2(_02081_),
    .ZN(_02082_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05596_ (.I0(\u_cpu.rf_ram.memory[104][5] ),
    .I1(\u_cpu.rf_ram.memory[105][5] ),
    .I2(\u_cpu.rf_ram.memory[106][5] ),
    .I3(\u_cpu.rf_ram.memory[107][5] ),
    .S0(_01615_),
    .S1(_01616_),
    .Z(_02083_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05597_ (.A1(_01594_),
    .A2(_02083_),
    .B(_01416_),
    .ZN(_02084_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05598_ (.I0(\u_cpu.rf_ram.memory[100][5] ),
    .I1(\u_cpu.rf_ram.memory[101][5] ),
    .I2(\u_cpu.rf_ram.memory[102][5] ),
    .I3(\u_cpu.rf_ram.memory[103][5] ),
    .S0(_01577_),
    .S1(_01549_),
    .Z(_02085_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05599_ (.A1(_01636_),
    .A2(_02085_),
    .ZN(_02086_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05600_ (.I0(\u_cpu.rf_ram.memory[96][5] ),
    .I1(\u_cpu.rf_ram.memory[97][5] ),
    .I2(\u_cpu.rf_ram.memory[98][5] ),
    .I3(\u_cpu.rf_ram.memory[99][5] ),
    .S0(_01602_),
    .S1(_01579_),
    .Z(_02087_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05601_ (.A1(_01594_),
    .A2(_02087_),
    .B(_01626_),
    .ZN(_02088_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _05602_ (.A1(_02082_),
    .A2(_02084_),
    .B1(_02086_),
    .B2(_02088_),
    .C(_01628_),
    .ZN(_02089_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05603_ (.I0(\u_cpu.rf_ram.memory[124][5] ),
    .I1(\u_cpu.rf_ram.memory[125][5] ),
    .I2(\u_cpu.rf_ram.memory[126][5] ),
    .I3(\u_cpu.rf_ram.memory[127][5] ),
    .S0(_01545_),
    .S1(_01642_),
    .Z(_02090_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05604_ (.A1(_01589_),
    .A2(_02090_),
    .ZN(_02091_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05605_ (.I0(\u_cpu.rf_ram.memory[120][5] ),
    .I1(\u_cpu.rf_ram.memory[121][5] ),
    .I2(\u_cpu.rf_ram.memory[122][5] ),
    .I3(\u_cpu.rf_ram.memory[123][5] ),
    .S0(_01646_),
    .S1(_01603_),
    .Z(_02092_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05606_ (.A1(_01601_),
    .A2(_02092_),
    .B(_01648_),
    .ZN(_02093_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05607_ (.I0(\u_cpu.rf_ram.memory[112][5] ),
    .I1(\u_cpu.rf_ram.memory[113][5] ),
    .I2(\u_cpu.rf_ram.memory[114][5] ),
    .I3(\u_cpu.rf_ram.memory[115][5] ),
    .S0(_01619_),
    .S1(_01620_),
    .Z(_02094_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05608_ (.A1(_01541_),
    .A2(_02094_),
    .ZN(_02095_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05609_ (.I0(\u_cpu.rf_ram.memory[116][5] ),
    .I1(\u_cpu.rf_ram.memory[117][5] ),
    .I2(\u_cpu.rf_ram.memory[118][5] ),
    .I3(\u_cpu.rf_ram.memory[119][5] ),
    .S0(_01623_),
    .S1(_01624_),
    .Z(_02096_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05610_ (.A1(_01614_),
    .A2(_02096_),
    .B(_01654_),
    .ZN(_02097_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _05611_ (.A1(_02091_),
    .A2(_02093_),
    .B1(_02095_),
    .B2(_02097_),
    .C(_01607_),
    .ZN(_02098_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _05612_ (.A1(_01422_),
    .A2(_02089_),
    .A3(_02098_),
    .ZN(_02099_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05613_ (.I0(\u_cpu.rf_ram.memory[92][5] ),
    .I1(\u_cpu.rf_ram.memory[93][5] ),
    .I2(\u_cpu.rf_ram.memory[94][5] ),
    .I3(\u_cpu.rf_ram.memory[95][5] ),
    .S0(_01610_),
    .S1(_01611_),
    .Z(_02100_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05614_ (.A1(_01398_),
    .A2(_02100_),
    .ZN(_02101_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05615_ (.I0(\u_cpu.rf_ram.memory[88][5] ),
    .I1(\u_cpu.rf_ram.memory[89][5] ),
    .I2(\u_cpu.rf_ram.memory[90][5] ),
    .I3(\u_cpu.rf_ram.memory[91][5] ),
    .S0(_01646_),
    .S1(_01603_),
    .Z(_02102_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05616_ (.A1(_01645_),
    .A2(_02102_),
    .B(_01648_),
    .ZN(_02103_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05617_ (.I0(\u_cpu.rf_ram.memory[80][5] ),
    .I1(\u_cpu.rf_ram.memory[81][5] ),
    .I2(\u_cpu.rf_ram.memory[82][5] ),
    .I3(\u_cpu.rf_ram.memory[83][5] ),
    .S0(_01590_),
    .S1(_01591_),
    .Z(_02104_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05618_ (.A1(_01609_),
    .A2(_02104_),
    .ZN(_02105_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05619_ (.I0(\u_cpu.rf_ram.memory[84][5] ),
    .I1(\u_cpu.rf_ram.memory[85][5] ),
    .I2(\u_cpu.rf_ram.memory[86][5] ),
    .I3(\u_cpu.rf_ram.memory[87][5] ),
    .S0(_01555_),
    .S1(_01652_),
    .Z(_02106_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05620_ (.A1(_01614_),
    .A2(_02106_),
    .B(_01654_),
    .ZN(_02107_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _05621_ (.A1(_02101_),
    .A2(_02103_),
    .B1(_02105_),
    .B2(_02107_),
    .C(_01426_),
    .ZN(_02108_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05622_ (.I0(\u_cpu.rf_ram.memory[64][5] ),
    .I1(\u_cpu.rf_ram.memory[65][5] ),
    .I2(\u_cpu.rf_ram.memory[66][5] ),
    .I3(\u_cpu.rf_ram.memory[67][5] ),
    .S0(_01571_),
    .S1(_01668_),
    .Z(_02109_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05623_ (.A1(_01667_),
    .A2(_02109_),
    .ZN(_02110_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05624_ (.I0(\u_cpu.rf_ram.memory[68][5] ),
    .I1(\u_cpu.rf_ram.memory[69][5] ),
    .I2(\u_cpu.rf_ram.memory[70][5] ),
    .I3(\u_cpu.rf_ram.memory[71][5] ),
    .S0(_01555_),
    .S1(_01652_),
    .Z(_02111_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05625_ (.A1(_01553_),
    .A2(_02111_),
    .B(_01565_),
    .ZN(_02112_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05626_ (.I0(\u_cpu.rf_ram.memory[72][5] ),
    .I1(\u_cpu.rf_ram.memory[73][5] ),
    .I2(\u_cpu.rf_ram.memory[74][5] ),
    .I3(\u_cpu.rf_ram.memory[75][5] ),
    .S0(_01610_),
    .S1(_01611_),
    .Z(_02113_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05627_ (.A1(_01667_),
    .A2(_02113_),
    .ZN(_02114_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05628_ (.I0(\u_cpu.rf_ram.memory[76][5] ),
    .I1(\u_cpu.rf_ram.memory[77][5] ),
    .I2(\u_cpu.rf_ram.memory[78][5] ),
    .I3(\u_cpu.rf_ram.memory[79][5] ),
    .S0(_01577_),
    .S1(_01549_),
    .Z(_02115_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05629_ (.A1(_01553_),
    .A2(_02115_),
    .B(_01417_),
    .ZN(_02116_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _05630_ (.A1(_02110_),
    .A2(_02112_),
    .B1(_02114_),
    .B2(_02116_),
    .C(_01568_),
    .ZN(_02117_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _05631_ (.A1(_01539_),
    .A2(_02108_),
    .A3(_02117_),
    .ZN(_02118_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05632_ (.A1(_02099_),
    .A2(_02118_),
    .B(_01402_),
    .ZN(_02119_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05633_ (.I0(\u_cpu.rf_ram.memory[136][5] ),
    .I1(\u_cpu.rf_ram.memory[137][5] ),
    .I2(\u_cpu.rf_ram.memory[138][5] ),
    .I3(\u_cpu.rf_ram.memory[139][5] ),
    .S0(_01680_),
    .S1(_01681_),
    .Z(_02120_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05634_ (.A1(_01399_),
    .A2(_02120_),
    .ZN(_02121_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05635_ (.I0(\u_cpu.rf_ram.memory[140][5] ),
    .I1(\u_cpu.rf_ram.memory[141][5] ),
    .I2(\u_cpu.rf_ram.memory[142][5] ),
    .I3(\u_cpu.rf_ram.memory[143][5] ),
    .S0(_01680_),
    .S1(_01681_),
    .Z(_02122_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05636_ (.A1(_01684_),
    .A2(_02122_),
    .B(_01582_),
    .ZN(_02123_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05637_ (.I0(\u_cpu.rf_ram.memory[128][5] ),
    .I1(\u_cpu.rf_ram.memory[129][5] ),
    .I2(\u_cpu.rf_ram.memory[130][5] ),
    .I3(\u_cpu.rf_ram.memory[131][5] ),
    .S0(_01687_),
    .S1(_01688_),
    .Z(_02124_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05638_ (.A1(_01399_),
    .A2(_02124_),
    .ZN(_02125_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05639_ (.I0(\u_cpu.rf_ram.memory[132][5] ),
    .I1(\u_cpu.rf_ram.memory[133][5] ),
    .I2(\u_cpu.rf_ram.memory[134][5] ),
    .I3(\u_cpu.rf_ram.memory[135][5] ),
    .S0(_01687_),
    .S1(_01688_),
    .Z(_02126_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05640_ (.A1(_01684_),
    .A2(_02126_),
    .B(_01418_),
    .ZN(_02127_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _05641_ (.A1(_02121_),
    .A2(_02123_),
    .B1(_02125_),
    .B2(_02127_),
    .C(_01404_),
    .ZN(_02128_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05642_ (.A1(_02119_),
    .A2(_02128_),
    .ZN(_02129_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05643_ (.A1(_01406_),
    .A2(_02080_),
    .B(_02129_),
    .ZN(_00005_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05644_ (.I0(\u_cpu.rf_ram.memory[8][6] ),
    .I1(\u_cpu.rf_ram.memory[9][6] ),
    .I2(\u_cpu.rf_ram.memory[10][6] ),
    .I3(\u_cpu.rf_ram.memory[11][6] ),
    .S0(_01546_),
    .S1(_01550_),
    .Z(_02130_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05645_ (.A1(_01542_),
    .A2(_02130_),
    .ZN(_02131_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05646_ (.I0(\u_cpu.rf_ram.memory[12][6] ),
    .I1(\u_cpu.rf_ram.memory[13][6] ),
    .I2(\u_cpu.rf_ram.memory[14][6] ),
    .I3(\u_cpu.rf_ram.memory[15][6] ),
    .S0(_01571_),
    .S1(_01557_),
    .Z(_02132_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05647_ (.A1(_01554_),
    .A2(_02132_),
    .B(_01417_),
    .ZN(_02133_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05648_ (.I0(\u_cpu.rf_ram.memory[4][6] ),
    .I1(\u_cpu.rf_ram.memory[5][6] ),
    .I2(\u_cpu.rf_ram.memory[6][6] ),
    .I3(\u_cpu.rf_ram.memory[7][6] ),
    .S0(_01578_),
    .S1(_01550_),
    .Z(_02134_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05649_ (.A1(_01554_),
    .A2(_02134_),
    .ZN(_02135_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05650_ (.I0(\u_cpu.rf_ram.memory[0][6] ),
    .I1(\u_cpu.rf_ram.memory[1][6] ),
    .I2(\u_cpu.rf_ram.memory[2][6] ),
    .I3(\u_cpu.rf_ram.memory[3][6] ),
    .S0(_01556_),
    .S1(_01557_),
    .Z(_02136_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05651_ (.A1(_01562_),
    .A2(_02136_),
    .B(_01565_),
    .ZN(_02137_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _05652_ (.A1(_02131_),
    .A2(_02133_),
    .B1(_02135_),
    .B2(_02137_),
    .C(_01568_),
    .ZN(_02138_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05653_ (.I0(\u_cpu.rf_ram.memory[20][6] ),
    .I1(\u_cpu.rf_ram.memory[21][6] ),
    .I2(\u_cpu.rf_ram.memory[22][6] ),
    .I3(\u_cpu.rf_ram.memory[23][6] ),
    .S0(_01572_),
    .S1(_01574_),
    .Z(_02139_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05654_ (.A1(_01570_),
    .A2(_02139_),
    .ZN(_02140_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05655_ (.I0(\u_cpu.rf_ram.memory[16][6] ),
    .I1(\u_cpu.rf_ram.memory[17][6] ),
    .I2(\u_cpu.rf_ram.memory[18][6] ),
    .I3(\u_cpu.rf_ram.memory[19][6] ),
    .S0(_01556_),
    .S1(_01580_),
    .Z(_02141_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05656_ (.A1(_01562_),
    .A2(_02141_),
    .B(_01582_),
    .ZN(_02142_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05657_ (.I0(\u_cpu.rf_ram.memory[28][6] ),
    .I1(\u_cpu.rf_ram.memory[29][6] ),
    .I2(\u_cpu.rf_ram.memory[30][6] ),
    .I3(\u_cpu.rf_ram.memory[31][6] ),
    .S0(_01546_),
    .S1(_01574_),
    .Z(_02143_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05658_ (.A1(_01570_),
    .A2(_02143_),
    .ZN(_02144_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05659_ (.I0(\u_cpu.rf_ram.memory[24][6] ),
    .I1(\u_cpu.rf_ram.memory[25][6] ),
    .I2(\u_cpu.rf_ram.memory[26][6] ),
    .I3(\u_cpu.rf_ram.memory[27][6] ),
    .S0(_01578_),
    .S1(_01580_),
    .Z(_02145_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05660_ (.A1(_01542_),
    .A2(_02145_),
    .B(_01418_),
    .ZN(_02146_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _05661_ (.A1(_02140_),
    .A2(_02142_),
    .B1(_02144_),
    .B2(_02146_),
    .C(_01426_),
    .ZN(_02147_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05662_ (.I0(\u_cpu.rf_ram.memory[52][6] ),
    .I1(\u_cpu.rf_ram.memory[53][6] ),
    .I2(\u_cpu.rf_ram.memory[54][6] ),
    .I3(\u_cpu.rf_ram.memory[55][6] ),
    .S0(_01590_),
    .S1(_01591_),
    .Z(_02148_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05663_ (.A1(_01589_),
    .A2(_02148_),
    .ZN(_02149_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05664_ (.I0(\u_cpu.rf_ram.memory[48][6] ),
    .I1(\u_cpu.rf_ram.memory[49][6] ),
    .I2(\u_cpu.rf_ram.memory[50][6] ),
    .I3(\u_cpu.rf_ram.memory[51][6] ),
    .S0(_01544_),
    .S1(_01548_),
    .Z(_02150_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05665_ (.A1(_01540_),
    .A2(_02150_),
    .B(_01564_),
    .ZN(_02151_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05666_ (.I0(\u_cpu.rf_ram.memory[60][6] ),
    .I1(\u_cpu.rf_ram.memory[61][6] ),
    .I2(\u_cpu.rf_ram.memory[62][6] ),
    .I3(\u_cpu.rf_ram.memory[63][6] ),
    .S0(_01598_),
    .S1(_01573_),
    .Z(_02152_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05667_ (.A1(_01636_),
    .A2(_02152_),
    .ZN(_02153_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05668_ (.I0(\u_cpu.rf_ram.memory[56][6] ),
    .I1(\u_cpu.rf_ram.memory[57][6] ),
    .I2(\u_cpu.rf_ram.memory[58][6] ),
    .I3(\u_cpu.rf_ram.memory[59][6] ),
    .S0(_01602_),
    .S1(_01579_),
    .Z(_02154_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05669_ (.A1(_01601_),
    .A2(_02154_),
    .B(_01605_),
    .ZN(_02155_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _05670_ (.A1(_02149_),
    .A2(_02151_),
    .B1(_02153_),
    .B2(_02155_),
    .C(_01607_),
    .ZN(_02156_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05671_ (.I0(\u_cpu.rf_ram.memory[40][6] ),
    .I1(\u_cpu.rf_ram.memory[41][6] ),
    .I2(\u_cpu.rf_ram.memory[42][6] ),
    .I3(\u_cpu.rf_ram.memory[43][6] ),
    .S0(_01545_),
    .S1(_01642_),
    .Z(_02157_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05672_ (.A1(_01609_),
    .A2(_02157_),
    .ZN(_02158_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05673_ (.I0(\u_cpu.rf_ram.memory[44][6] ),
    .I1(\u_cpu.rf_ram.memory[45][6] ),
    .I2(\u_cpu.rf_ram.memory[46][6] ),
    .I3(\u_cpu.rf_ram.memory[47][6] ),
    .S0(_01615_),
    .S1(_01616_),
    .Z(_02159_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05674_ (.A1(_01397_),
    .A2(_02159_),
    .B(_01416_),
    .ZN(_02160_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05675_ (.I0(\u_cpu.rf_ram.memory[36][6] ),
    .I1(\u_cpu.rf_ram.memory[37][6] ),
    .I2(\u_cpu.rf_ram.memory[38][6] ),
    .I3(\u_cpu.rf_ram.memory[39][6] ),
    .S0(_01619_),
    .S1(_01620_),
    .Z(_02161_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05676_ (.A1(_01597_),
    .A2(_02161_),
    .ZN(_02162_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05677_ (.I0(\u_cpu.rf_ram.memory[32][6] ),
    .I1(\u_cpu.rf_ram.memory[33][6] ),
    .I2(\u_cpu.rf_ram.memory[34][6] ),
    .I3(\u_cpu.rf_ram.memory[35][6] ),
    .S0(_01623_),
    .S1(_01624_),
    .Z(_02163_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05678_ (.A1(_01645_),
    .A2(_02163_),
    .B(_01626_),
    .ZN(_02164_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _05679_ (.A1(_02158_),
    .A2(_02160_),
    .B1(_02162_),
    .B2(_02164_),
    .C(_01628_),
    .ZN(_02165_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _05680_ (.A1(_01422_),
    .A2(_02156_),
    .A3(_02165_),
    .Z(_02166_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _05681_ (.A1(_01539_),
    .A2(_02138_),
    .A3(_02147_),
    .B(_02166_),
    .ZN(_02167_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05682_ (.I0(\u_cpu.rf_ram.memory[108][6] ),
    .I1(\u_cpu.rf_ram.memory[109][6] ),
    .I2(\u_cpu.rf_ram.memory[110][6] ),
    .I3(\u_cpu.rf_ram.memory[111][6] ),
    .S0(_01598_),
    .S1(_01573_),
    .Z(_02168_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05683_ (.A1(_01597_),
    .A2(_02168_),
    .ZN(_02169_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05684_ (.I0(\u_cpu.rf_ram.memory[104][6] ),
    .I1(\u_cpu.rf_ram.memory[105][6] ),
    .I2(\u_cpu.rf_ram.memory[106][6] ),
    .I3(\u_cpu.rf_ram.memory[107][6] ),
    .S0(_01615_),
    .S1(_01616_),
    .Z(_02170_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05685_ (.A1(_01594_),
    .A2(_02170_),
    .B(_01416_),
    .ZN(_02171_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05686_ (.I0(\u_cpu.rf_ram.memory[100][6] ),
    .I1(\u_cpu.rf_ram.memory[101][6] ),
    .I2(\u_cpu.rf_ram.memory[102][6] ),
    .I3(\u_cpu.rf_ram.memory[103][6] ),
    .S0(_01577_),
    .S1(_01549_),
    .Z(_02172_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05687_ (.A1(_01636_),
    .A2(_02172_),
    .ZN(_02173_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05688_ (.I0(\u_cpu.rf_ram.memory[96][6] ),
    .I1(\u_cpu.rf_ram.memory[97][6] ),
    .I2(\u_cpu.rf_ram.memory[98][6] ),
    .I3(\u_cpu.rf_ram.memory[99][6] ),
    .S0(_01602_),
    .S1(_01579_),
    .Z(_02174_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05689_ (.A1(_01594_),
    .A2(_02174_),
    .B(_01626_),
    .ZN(_02175_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _05690_ (.A1(_02169_),
    .A2(_02171_),
    .B1(_02173_),
    .B2(_02175_),
    .C(_01628_),
    .ZN(_02176_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05691_ (.I0(\u_cpu.rf_ram.memory[124][6] ),
    .I1(\u_cpu.rf_ram.memory[125][6] ),
    .I2(\u_cpu.rf_ram.memory[126][6] ),
    .I3(\u_cpu.rf_ram.memory[127][6] ),
    .S0(_01545_),
    .S1(_01642_),
    .Z(_02177_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05692_ (.A1(_01589_),
    .A2(_02177_),
    .ZN(_02178_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05693_ (.I0(\u_cpu.rf_ram.memory[120][6] ),
    .I1(\u_cpu.rf_ram.memory[121][6] ),
    .I2(\u_cpu.rf_ram.memory[122][6] ),
    .I3(\u_cpu.rf_ram.memory[123][6] ),
    .S0(_01646_),
    .S1(_01603_),
    .Z(_02179_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05694_ (.A1(_01601_),
    .A2(_02179_),
    .B(_01605_),
    .ZN(_02180_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05695_ (.I0(\u_cpu.rf_ram.memory[112][6] ),
    .I1(\u_cpu.rf_ram.memory[113][6] ),
    .I2(\u_cpu.rf_ram.memory[114][6] ),
    .I3(\u_cpu.rf_ram.memory[115][6] ),
    .S0(_01619_),
    .S1(_01620_),
    .Z(_02181_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05696_ (.A1(_01541_),
    .A2(_02181_),
    .ZN(_02182_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05697_ (.I0(\u_cpu.rf_ram.memory[116][6] ),
    .I1(\u_cpu.rf_ram.memory[117][6] ),
    .I2(\u_cpu.rf_ram.memory[118][6] ),
    .I3(\u_cpu.rf_ram.memory[119][6] ),
    .S0(_01623_),
    .S1(_01624_),
    .Z(_02183_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05698_ (.A1(_01614_),
    .A2(_02183_),
    .B(_01654_),
    .ZN(_02184_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _05699_ (.A1(_02178_),
    .A2(_02180_),
    .B1(_02182_),
    .B2(_02184_),
    .C(_01607_),
    .ZN(_02185_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _05700_ (.A1(_01422_),
    .A2(_02176_),
    .A3(_02185_),
    .ZN(_02186_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05701_ (.I0(\u_cpu.rf_ram.memory[92][6] ),
    .I1(\u_cpu.rf_ram.memory[93][6] ),
    .I2(\u_cpu.rf_ram.memory[94][6] ),
    .I3(\u_cpu.rf_ram.memory[95][6] ),
    .S0(_01610_),
    .S1(_01611_),
    .Z(_02187_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05702_ (.A1(_01398_),
    .A2(_02187_),
    .ZN(_02188_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05703_ (.I0(\u_cpu.rf_ram.memory[88][6] ),
    .I1(\u_cpu.rf_ram.memory[89][6] ),
    .I2(\u_cpu.rf_ram.memory[90][6] ),
    .I3(\u_cpu.rf_ram.memory[91][6] ),
    .S0(_01646_),
    .S1(_01603_),
    .Z(_02189_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05704_ (.A1(_01645_),
    .A2(_02189_),
    .B(_01648_),
    .ZN(_02190_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05705_ (.I0(\u_cpu.rf_ram.memory[80][6] ),
    .I1(\u_cpu.rf_ram.memory[81][6] ),
    .I2(\u_cpu.rf_ram.memory[82][6] ),
    .I3(\u_cpu.rf_ram.memory[83][6] ),
    .S0(_01590_),
    .S1(_01591_),
    .Z(_02191_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05706_ (.A1(_01609_),
    .A2(_02191_),
    .ZN(_02192_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05707_ (.I0(\u_cpu.rf_ram.memory[84][6] ),
    .I1(\u_cpu.rf_ram.memory[85][6] ),
    .I2(\u_cpu.rf_ram.memory[86][6] ),
    .I3(\u_cpu.rf_ram.memory[87][6] ),
    .S0(_01555_),
    .S1(_01652_),
    .Z(_02193_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05708_ (.A1(_01614_),
    .A2(_02193_),
    .B(_01654_),
    .ZN(_02194_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _05709_ (.A1(_02188_),
    .A2(_02190_),
    .B1(_02192_),
    .B2(_02194_),
    .C(_01426_),
    .ZN(_02195_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05710_ (.I0(\u_cpu.rf_ram.memory[64][6] ),
    .I1(\u_cpu.rf_ram.memory[65][6] ),
    .I2(\u_cpu.rf_ram.memory[66][6] ),
    .I3(\u_cpu.rf_ram.memory[67][6] ),
    .S0(_01571_),
    .S1(_01668_),
    .Z(_02196_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05711_ (.A1(_01667_),
    .A2(_02196_),
    .ZN(_02197_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05712_ (.I0(\u_cpu.rf_ram.memory[68][6] ),
    .I1(\u_cpu.rf_ram.memory[69][6] ),
    .I2(\u_cpu.rf_ram.memory[70][6] ),
    .I3(\u_cpu.rf_ram.memory[71][6] ),
    .S0(_01555_),
    .S1(_01652_),
    .Z(_02198_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05713_ (.A1(_01553_),
    .A2(_02198_),
    .B(_01565_),
    .ZN(_02199_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05714_ (.I0(\u_cpu.rf_ram.memory[72][6] ),
    .I1(\u_cpu.rf_ram.memory[73][6] ),
    .I2(\u_cpu.rf_ram.memory[74][6] ),
    .I3(\u_cpu.rf_ram.memory[75][6] ),
    .S0(_01610_),
    .S1(_01611_),
    .Z(_02200_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05715_ (.A1(_01667_),
    .A2(_02200_),
    .ZN(_02201_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05716_ (.I0(\u_cpu.rf_ram.memory[76][6] ),
    .I1(\u_cpu.rf_ram.memory[77][6] ),
    .I2(\u_cpu.rf_ram.memory[78][6] ),
    .I3(\u_cpu.rf_ram.memory[79][6] ),
    .S0(_01577_),
    .S1(_01549_),
    .Z(_02202_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05717_ (.A1(_01553_),
    .A2(_02202_),
    .B(_01648_),
    .ZN(_02203_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _05718_ (.A1(_02197_),
    .A2(_02199_),
    .B1(_02201_),
    .B2(_02203_),
    .C(_01568_),
    .ZN(_02204_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _05719_ (.A1(_01539_),
    .A2(_02195_),
    .A3(_02204_),
    .ZN(_02205_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05720_ (.A1(_02186_),
    .A2(_02205_),
    .B(_01402_),
    .ZN(_02206_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05721_ (.I0(\u_cpu.rf_ram.memory[136][6] ),
    .I1(\u_cpu.rf_ram.memory[137][6] ),
    .I2(\u_cpu.rf_ram.memory[138][6] ),
    .I3(\u_cpu.rf_ram.memory[139][6] ),
    .S0(_01687_),
    .S1(_01681_),
    .Z(_02207_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05722_ (.A1(_01399_),
    .A2(_02207_),
    .ZN(_02208_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05723_ (.I0(\u_cpu.rf_ram.memory[140][6] ),
    .I1(\u_cpu.rf_ram.memory[141][6] ),
    .I2(\u_cpu.rf_ram.memory[142][6] ),
    .I3(\u_cpu.rf_ram.memory[143][6] ),
    .S0(_01680_),
    .S1(_01681_),
    .Z(_02209_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05724_ (.A1(_01684_),
    .A2(_02209_),
    .B(_01582_),
    .ZN(_02210_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05725_ (.I0(\u_cpu.rf_ram.memory[128][6] ),
    .I1(\u_cpu.rf_ram.memory[129][6] ),
    .I2(\u_cpu.rf_ram.memory[130][6] ),
    .I3(\u_cpu.rf_ram.memory[131][6] ),
    .S0(_01572_),
    .S1(_01688_),
    .Z(_02211_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05726_ (.A1(_01399_),
    .A2(_02211_),
    .ZN(_02212_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05727_ (.I0(\u_cpu.rf_ram.memory[132][6] ),
    .I1(\u_cpu.rf_ram.memory[133][6] ),
    .I2(\u_cpu.rf_ram.memory[134][6] ),
    .I3(\u_cpu.rf_ram.memory[135][6] ),
    .S0(_01687_),
    .S1(_01688_),
    .Z(_02213_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05728_ (.A1(_01684_),
    .A2(_02213_),
    .B(_01418_),
    .ZN(_02214_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _05729_ (.A1(_02208_),
    .A2(_02210_),
    .B1(_02212_),
    .B2(_02214_),
    .C(_01404_),
    .ZN(_02215_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05730_ (.A1(_02206_),
    .A2(_02215_),
    .ZN(_02216_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05731_ (.A1(_01406_),
    .A2(_02167_),
    .B(_02216_),
    .ZN(_00006_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05732_ (.I0(\u_cpu.rf_ram.memory[8][7] ),
    .I1(\u_cpu.rf_ram.memory[9][7] ),
    .I2(\u_cpu.rf_ram.memory[10][7] ),
    .I3(\u_cpu.rf_ram.memory[11][7] ),
    .S0(_01546_),
    .S1(_01550_),
    .Z(_02217_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05733_ (.A1(_01542_),
    .A2(_02217_),
    .ZN(_02218_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05734_ (.I0(\u_cpu.rf_ram.memory[12][7] ),
    .I1(\u_cpu.rf_ram.memory[13][7] ),
    .I2(\u_cpu.rf_ram.memory[14][7] ),
    .I3(\u_cpu.rf_ram.memory[15][7] ),
    .S0(_01571_),
    .S1(_01668_),
    .Z(_02219_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05735_ (.A1(_01398_),
    .A2(_02219_),
    .B(_01417_),
    .ZN(_02220_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05736_ (.I0(\u_cpu.rf_ram.memory[4][7] ),
    .I1(\u_cpu.rf_ram.memory[5][7] ),
    .I2(\u_cpu.rf_ram.memory[6][7] ),
    .I3(\u_cpu.rf_ram.memory[7][7] ),
    .S0(_01578_),
    .S1(_01580_),
    .Z(_02221_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05737_ (.A1(_01554_),
    .A2(_02221_),
    .ZN(_02222_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05738_ (.I0(\u_cpu.rf_ram.memory[0][7] ),
    .I1(\u_cpu.rf_ram.memory[1][7] ),
    .I2(\u_cpu.rf_ram.memory[2][7] ),
    .I3(\u_cpu.rf_ram.memory[3][7] ),
    .S0(_01556_),
    .S1(_01557_),
    .Z(_02223_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05739_ (.A1(_01562_),
    .A2(_02223_),
    .B(_01565_),
    .ZN(_02224_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _05740_ (.A1(_02218_),
    .A2(_02220_),
    .B1(_02222_),
    .B2(_02224_),
    .C(_01568_),
    .ZN(_02225_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05741_ (.I0(\u_cpu.rf_ram.memory[20][7] ),
    .I1(\u_cpu.rf_ram.memory[21][7] ),
    .I2(\u_cpu.rf_ram.memory[22][7] ),
    .I3(\u_cpu.rf_ram.memory[23][7] ),
    .S0(_01572_),
    .S1(_01574_),
    .Z(_02226_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05742_ (.A1(_01570_),
    .A2(_02226_),
    .ZN(_02227_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05743_ (.I0(\u_cpu.rf_ram.memory[16][7] ),
    .I1(\u_cpu.rf_ram.memory[17][7] ),
    .I2(\u_cpu.rf_ram.memory[18][7] ),
    .I3(\u_cpu.rf_ram.memory[19][7] ),
    .S0(_01556_),
    .S1(_01557_),
    .Z(_02228_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05744_ (.A1(_01562_),
    .A2(_02228_),
    .B(_01582_),
    .ZN(_02229_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05745_ (.I0(\u_cpu.rf_ram.memory[28][7] ),
    .I1(\u_cpu.rf_ram.memory[29][7] ),
    .I2(\u_cpu.rf_ram.memory[30][7] ),
    .I3(\u_cpu.rf_ram.memory[31][7] ),
    .S0(_01546_),
    .S1(_01550_),
    .Z(_02230_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05746_ (.A1(_01554_),
    .A2(_02230_),
    .ZN(_02231_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05747_ (.I0(\u_cpu.rf_ram.memory[24][7] ),
    .I1(\u_cpu.rf_ram.memory[25][7] ),
    .I2(\u_cpu.rf_ram.memory[26][7] ),
    .I3(\u_cpu.rf_ram.memory[27][7] ),
    .S0(_01578_),
    .S1(_01580_),
    .Z(_02232_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05748_ (.A1(_01542_),
    .A2(_02232_),
    .B(_01417_),
    .ZN(_02233_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _05749_ (.A1(_02227_),
    .A2(_02229_),
    .B1(_02231_),
    .B2(_02233_),
    .C(_01426_),
    .ZN(_02234_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05750_ (.I0(\u_cpu.rf_ram.memory[52][7] ),
    .I1(\u_cpu.rf_ram.memory[53][7] ),
    .I2(\u_cpu.rf_ram.memory[54][7] ),
    .I3(\u_cpu.rf_ram.memory[55][7] ),
    .S0(_01590_),
    .S1(_01591_),
    .Z(_02235_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05751_ (.A1(_01589_),
    .A2(_02235_),
    .ZN(_02236_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05752_ (.I0(\u_cpu.rf_ram.memory[48][7] ),
    .I1(\u_cpu.rf_ram.memory[49][7] ),
    .I2(\u_cpu.rf_ram.memory[50][7] ),
    .I3(\u_cpu.rf_ram.memory[51][7] ),
    .S0(_01544_),
    .S1(_01548_),
    .Z(_02237_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05753_ (.A1(_01540_),
    .A2(_02237_),
    .B(_01564_),
    .ZN(_02238_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05754_ (.I0(\u_cpu.rf_ram.memory[60][7] ),
    .I1(\u_cpu.rf_ram.memory[61][7] ),
    .I2(\u_cpu.rf_ram.memory[62][7] ),
    .I3(\u_cpu.rf_ram.memory[63][7] ),
    .S0(_01598_),
    .S1(_01573_),
    .Z(_02239_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05755_ (.A1(_01636_),
    .A2(_02239_),
    .ZN(_02240_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05756_ (.I0(\u_cpu.rf_ram.memory[56][7] ),
    .I1(\u_cpu.rf_ram.memory[57][7] ),
    .I2(\u_cpu.rf_ram.memory[58][7] ),
    .I3(\u_cpu.rf_ram.memory[59][7] ),
    .S0(_01602_),
    .S1(_01579_),
    .Z(_02241_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05757_ (.A1(_01601_),
    .A2(_02241_),
    .B(_01605_),
    .ZN(_02242_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _05758_ (.A1(_02236_),
    .A2(_02238_),
    .B1(_02240_),
    .B2(_02242_),
    .C(_01425_),
    .ZN(_02243_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05759_ (.I0(\u_cpu.rf_ram.memory[40][7] ),
    .I1(\u_cpu.rf_ram.memory[41][7] ),
    .I2(\u_cpu.rf_ram.memory[42][7] ),
    .I3(\u_cpu.rf_ram.memory[43][7] ),
    .S0(_01545_),
    .S1(_01642_),
    .Z(_02244_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05760_ (.A1(_01609_),
    .A2(_02244_),
    .ZN(_02245_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05761_ (.I0(\u_cpu.rf_ram.memory[44][7] ),
    .I1(\u_cpu.rf_ram.memory[45][7] ),
    .I2(\u_cpu.rf_ram.memory[46][7] ),
    .I3(\u_cpu.rf_ram.memory[47][7] ),
    .S0(_01615_),
    .S1(_01616_),
    .Z(_02246_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05762_ (.A1(_01397_),
    .A2(_02246_),
    .B(_01416_),
    .ZN(_02247_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05763_ (.I0(\u_cpu.rf_ram.memory[36][7] ),
    .I1(\u_cpu.rf_ram.memory[37][7] ),
    .I2(\u_cpu.rf_ram.memory[38][7] ),
    .I3(\u_cpu.rf_ram.memory[39][7] ),
    .S0(_01619_),
    .S1(_01620_),
    .Z(_02248_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05764_ (.A1(_01597_),
    .A2(_02248_),
    .ZN(_02249_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05765_ (.I0(\u_cpu.rf_ram.memory[32][7] ),
    .I1(\u_cpu.rf_ram.memory[33][7] ),
    .I2(\u_cpu.rf_ram.memory[34][7] ),
    .I3(\u_cpu.rf_ram.memory[35][7] ),
    .S0(_01623_),
    .S1(_01624_),
    .Z(_02250_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05766_ (.A1(_01645_),
    .A2(_02250_),
    .B(_01626_),
    .ZN(_02251_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _05767_ (.A1(_02245_),
    .A2(_02247_),
    .B1(_02249_),
    .B2(_02251_),
    .C(_01628_),
    .ZN(_02252_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _05768_ (.A1(_01421_),
    .A2(_02243_),
    .A3(_02252_),
    .Z(_02253_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _05769_ (.A1(_01539_),
    .A2(_02225_),
    .A3(_02234_),
    .B(_02253_),
    .ZN(_02254_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05770_ (.I0(\u_cpu.rf_ram.memory[108][7] ),
    .I1(\u_cpu.rf_ram.memory[109][7] ),
    .I2(\u_cpu.rf_ram.memory[110][7] ),
    .I3(\u_cpu.rf_ram.memory[111][7] ),
    .S0(_01598_),
    .S1(_01573_),
    .Z(_02255_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05771_ (.A1(_01597_),
    .A2(_02255_),
    .ZN(_02256_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05772_ (.I0(\u_cpu.rf_ram.memory[104][7] ),
    .I1(\u_cpu.rf_ram.memory[105][7] ),
    .I2(\u_cpu.rf_ram.memory[106][7] ),
    .I3(\u_cpu.rf_ram.memory[107][7] ),
    .S0(_01615_),
    .S1(_01616_),
    .Z(_02257_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05773_ (.A1(_01594_),
    .A2(_02257_),
    .B(_01416_),
    .ZN(_02258_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05774_ (.I0(\u_cpu.rf_ram.memory[100][7] ),
    .I1(\u_cpu.rf_ram.memory[101][7] ),
    .I2(\u_cpu.rf_ram.memory[102][7] ),
    .I3(\u_cpu.rf_ram.memory[103][7] ),
    .S0(_01577_),
    .S1(_01549_),
    .Z(_02259_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05775_ (.A1(_01636_),
    .A2(_02259_),
    .ZN(_02260_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05776_ (.I0(\u_cpu.rf_ram.memory[96][7] ),
    .I1(\u_cpu.rf_ram.memory[97][7] ),
    .I2(\u_cpu.rf_ram.memory[98][7] ),
    .I3(\u_cpu.rf_ram.memory[99][7] ),
    .S0(_01602_),
    .S1(_01579_),
    .Z(_02261_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05777_ (.A1(_01594_),
    .A2(_02261_),
    .B(_01564_),
    .ZN(_02262_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _05778_ (.A1(_02256_),
    .A2(_02258_),
    .B1(_02260_),
    .B2(_02262_),
    .C(_01628_),
    .ZN(_02263_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05779_ (.I0(\u_cpu.rf_ram.memory[124][7] ),
    .I1(\u_cpu.rf_ram.memory[125][7] ),
    .I2(\u_cpu.rf_ram.memory[126][7] ),
    .I3(\u_cpu.rf_ram.memory[127][7] ),
    .S0(_01545_),
    .S1(_01642_),
    .Z(_02264_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05780_ (.A1(_01589_),
    .A2(_02264_),
    .ZN(_02265_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05781_ (.I0(\u_cpu.rf_ram.memory[120][7] ),
    .I1(\u_cpu.rf_ram.memory[121][7] ),
    .I2(\u_cpu.rf_ram.memory[122][7] ),
    .I3(\u_cpu.rf_ram.memory[123][7] ),
    .S0(_01646_),
    .S1(_01603_),
    .Z(_02266_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05782_ (.A1(_01601_),
    .A2(_02266_),
    .B(_01605_),
    .ZN(_02267_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05783_ (.I0(\u_cpu.rf_ram.memory[112][7] ),
    .I1(\u_cpu.rf_ram.memory[113][7] ),
    .I2(\u_cpu.rf_ram.memory[114][7] ),
    .I3(\u_cpu.rf_ram.memory[115][7] ),
    .S0(_01619_),
    .S1(_01620_),
    .Z(_02268_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05784_ (.A1(_01541_),
    .A2(_02268_),
    .ZN(_02269_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05785_ (.I0(\u_cpu.rf_ram.memory[116][7] ),
    .I1(\u_cpu.rf_ram.memory[117][7] ),
    .I2(\u_cpu.rf_ram.memory[118][7] ),
    .I3(\u_cpu.rf_ram.memory[119][7] ),
    .S0(_01623_),
    .S1(_01624_),
    .Z(_02270_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05786_ (.A1(_01614_),
    .A2(_02270_),
    .B(_01626_),
    .ZN(_02271_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _05787_ (.A1(_02265_),
    .A2(_02267_),
    .B1(_02269_),
    .B2(_02271_),
    .C(_01607_),
    .ZN(_02272_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _05788_ (.A1(_01422_),
    .A2(_02263_),
    .A3(_02272_),
    .ZN(_02273_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05789_ (.I0(\u_cpu.rf_ram.memory[92][7] ),
    .I1(\u_cpu.rf_ram.memory[93][7] ),
    .I2(\u_cpu.rf_ram.memory[94][7] ),
    .I3(\u_cpu.rf_ram.memory[95][7] ),
    .S0(_01610_),
    .S1(_01611_),
    .Z(_02274_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05790_ (.A1(_01398_),
    .A2(_02274_),
    .ZN(_02275_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05791_ (.I0(\u_cpu.rf_ram.memory[88][7] ),
    .I1(\u_cpu.rf_ram.memory[89][7] ),
    .I2(\u_cpu.rf_ram.memory[90][7] ),
    .I3(\u_cpu.rf_ram.memory[91][7] ),
    .S0(_01646_),
    .S1(_01603_),
    .Z(_02276_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05792_ (.A1(_01645_),
    .A2(_02276_),
    .B(_01648_),
    .ZN(_02277_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05793_ (.I0(\u_cpu.rf_ram.memory[80][7] ),
    .I1(\u_cpu.rf_ram.memory[81][7] ),
    .I2(\u_cpu.rf_ram.memory[82][7] ),
    .I3(\u_cpu.rf_ram.memory[83][7] ),
    .S0(_01590_),
    .S1(_01591_),
    .Z(_02278_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05794_ (.A1(_01541_),
    .A2(_02278_),
    .ZN(_02279_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05795_ (.I0(\u_cpu.rf_ram.memory[84][7] ),
    .I1(\u_cpu.rf_ram.memory[85][7] ),
    .I2(\u_cpu.rf_ram.memory[86][7] ),
    .I3(\u_cpu.rf_ram.memory[87][7] ),
    .S0(_01555_),
    .S1(_01652_),
    .Z(_02280_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05796_ (.A1(_01614_),
    .A2(_02280_),
    .B(_01654_),
    .ZN(_02281_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _05797_ (.A1(_02275_),
    .A2(_02277_),
    .B1(_02279_),
    .B2(_02281_),
    .C(_01607_),
    .ZN(_02282_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05798_ (.I0(\u_cpu.rf_ram.memory[64][7] ),
    .I1(\u_cpu.rf_ram.memory[65][7] ),
    .I2(\u_cpu.rf_ram.memory[66][7] ),
    .I3(\u_cpu.rf_ram.memory[67][7] ),
    .S0(_01571_),
    .S1(_01668_),
    .Z(_02283_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05799_ (.A1(_01667_),
    .A2(_02283_),
    .ZN(_02284_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05800_ (.I0(\u_cpu.rf_ram.memory[68][7] ),
    .I1(\u_cpu.rf_ram.memory[69][7] ),
    .I2(\u_cpu.rf_ram.memory[70][7] ),
    .I3(\u_cpu.rf_ram.memory[71][7] ),
    .S0(_01555_),
    .S1(_01652_),
    .Z(_02285_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05801_ (.A1(_01553_),
    .A2(_02285_),
    .B(_01654_),
    .ZN(_02286_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05802_ (.I0(\u_cpu.rf_ram.memory[72][7] ),
    .I1(\u_cpu.rf_ram.memory[73][7] ),
    .I2(\u_cpu.rf_ram.memory[74][7] ),
    .I3(\u_cpu.rf_ram.memory[75][7] ),
    .S0(_01610_),
    .S1(_01611_),
    .Z(_02287_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05803_ (.A1(_01609_),
    .A2(_02287_),
    .ZN(_02288_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05804_ (.I0(\u_cpu.rf_ram.memory[76][7] ),
    .I1(\u_cpu.rf_ram.memory[77][7] ),
    .I2(\u_cpu.rf_ram.memory[78][7] ),
    .I3(\u_cpu.rf_ram.memory[79][7] ),
    .S0(_01577_),
    .S1(_01549_),
    .Z(_02289_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05805_ (.A1(_01553_),
    .A2(_02289_),
    .B(_01648_),
    .ZN(_02290_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _05806_ (.A1(_02284_),
    .A2(_02286_),
    .B1(_02288_),
    .B2(_02290_),
    .C(_01568_),
    .ZN(_02291_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _05807_ (.A1(_01539_),
    .A2(_02282_),
    .A3(_02291_),
    .ZN(_02292_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05808_ (.A1(_02273_),
    .A2(_02292_),
    .B(_01402_),
    .ZN(_02293_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05809_ (.I0(\u_cpu.rf_ram.memory[136][7] ),
    .I1(\u_cpu.rf_ram.memory[137][7] ),
    .I2(\u_cpu.rf_ram.memory[138][7] ),
    .I3(\u_cpu.rf_ram.memory[139][7] ),
    .S0(_01687_),
    .S1(_01688_),
    .Z(_02294_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05810_ (.A1(_01399_),
    .A2(_02294_),
    .ZN(_02295_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05811_ (.I0(\u_cpu.rf_ram.memory[140][7] ),
    .I1(\u_cpu.rf_ram.memory[141][7] ),
    .I2(\u_cpu.rf_ram.memory[142][7] ),
    .I3(\u_cpu.rf_ram.memory[143][7] ),
    .S0(_01680_),
    .S1(_01681_),
    .Z(_02296_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05812_ (.A1(_01684_),
    .A2(_02296_),
    .B(_01582_),
    .ZN(_02297_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05813_ (.I0(\u_cpu.rf_ram.memory[128][7] ),
    .I1(\u_cpu.rf_ram.memory[129][7] ),
    .I2(\u_cpu.rf_ram.memory[130][7] ),
    .I3(\u_cpu.rf_ram.memory[131][7] ),
    .S0(_01572_),
    .S1(_01574_),
    .Z(_02298_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05814_ (.A1(_01570_),
    .A2(_02298_),
    .ZN(_02299_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05815_ (.I0(\u_cpu.rf_ram.memory[132][7] ),
    .I1(\u_cpu.rf_ram.memory[133][7] ),
    .I2(\u_cpu.rf_ram.memory[134][7] ),
    .I3(\u_cpu.rf_ram.memory[135][7] ),
    .S0(_01687_),
    .S1(_01688_),
    .Z(_02300_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05816_ (.A1(_01684_),
    .A2(_02300_),
    .B(_01418_),
    .ZN(_02301_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _05817_ (.A1(_02295_),
    .A2(_02297_),
    .B1(_02299_),
    .B2(_02301_),
    .C(_01404_),
    .ZN(_02302_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05818_ (.A1(_02293_),
    .A2(_02302_),
    .ZN(_02303_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05819_ (.A1(_01406_),
    .A2(_02254_),
    .B(_02303_),
    .ZN(_00007_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _05820_ (.A1(\u_cpu.cpu.state.o_cnt_r[0] ),
    .A2(\u_cpu.cpu.state.o_cnt_r[1] ),
    .A3(\u_cpu.cpu.state.o_cnt_r[2] ),
    .A4(\u_cpu.cpu.state.o_cnt_r[3] ),
    .Z(_02304_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05821_ (.I(_02304_),
    .Z(_02305_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05822_ (.I(\u_arbiter.i_wb_cpu_dbus_we ),
    .Z(_02306_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05823_ (.I(_01409_),
    .ZN(_02307_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _05824_ (.A1(_02306_),
    .A2(\u_cpu.cpu.bufreg.i_sh_signed ),
    .B(_02307_),
    .C(_01374_),
    .ZN(_02308_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05825_ (.I(\u_cpu.cpu.alu.i_rs1 ),
    .Z(_02309_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05826_ (.A1(_02309_),
    .A2(\u_cpu.cpu.alu.add_cy_r ),
    .ZN(_02310_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05827_ (.I(\u_cpu.cpu.bufreg2.i_cnt_done ),
    .Z(_02311_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05828_ (.I(\u_cpu.cpu.immdec.imm11_7[0] ),
    .ZN(_02312_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05829_ (.I(\u_cpu.cpu.decode.opcode[0] ),
    .Z(_02313_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _05830_ (.A1(_01372_),
    .A2(\u_cpu.cpu.decode.opcode[1] ),
    .A3(_02313_),
    .ZN(_02314_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _05831_ (.A1(_02306_),
    .A2(_02312_),
    .A3(_02314_),
    .Z(_02315_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05832_ (.A1(_02306_),
    .A2(_02314_),
    .B(\u_cpu.cpu.immdec.imm24_20[0] ),
    .ZN(_02316_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _05833_ (.A1(_01369_),
    .A2(_01372_),
    .A3(_01374_),
    .ZN(_02317_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _05834_ (.A1(_02311_),
    .A2(\u_cpu.cpu.immdec.imm31 ),
    .A3(_02317_),
    .ZN(_02318_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _05835_ (.A1(_02311_),
    .A2(_02315_),
    .A3(_02316_),
    .B(_02318_),
    .ZN(_02319_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05836_ (.I(\u_cpu.rf_ram_if.rtrig1 ),
    .Z(_02320_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _05837_ (.I(\u_cpu.rf_ram.regzero ),
    .ZN(_02321_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05838_ (.A1(\u_cpu.rf_ram.rdata[0] ),
    .A2(_02321_),
    .ZN(_02322_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05839_ (.A1(\u_cpu.rf_ram_if.rdata1[0] ),
    .A2(_02320_),
    .ZN(_02323_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05840_ (.A1(_02320_),
    .A2(_02322_),
    .B(_02323_),
    .ZN(_02324_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05841_ (.I0(_02319_),
    .I1(_02324_),
    .S(_02306_),
    .Z(_02325_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _05842_ (.A1(_02308_),
    .A2(_02325_),
    .Z(_02326_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05843_ (.A1(_02309_),
    .A2(\u_cpu.cpu.alu.add_cy_r ),
    .ZN(_02327_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05844_ (.A1(_02310_),
    .A2(_02326_),
    .B(_02327_),
    .ZN(_02328_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05845_ (.A1(_02305_),
    .A2(_02328_),
    .ZN(_02329_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05846_ (.A1(_02305_),
    .A2(_02308_),
    .B(_02329_),
    .ZN(_00021_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05847_ (.A1(_01369_),
    .A2(_01390_),
    .ZN(_02330_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05848_ (.A1(_01369_),
    .A2(_02309_),
    .B(_02330_),
    .ZN(_02331_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _05849_ (.I(_01370_),
    .ZN(_02332_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05850_ (.I(\u_cpu.cpu.bne_or_bge ),
    .ZN(_02333_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05851_ (.A1(_02332_),
    .A2(_02333_),
    .ZN(_02334_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05852_ (.A1(_01370_),
    .A2(_02331_),
    .B(_02333_),
    .ZN(_02335_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _05853_ (.A1(_01379_),
    .A2(_01382_),
    .Z(_02336_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05854_ (.I(\u_cpu.cpu.decode.op22 ),
    .ZN(_02337_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _05855_ (.A1(\u_cpu.cpu.mem_bytecnt[1] ),
    .A2(\u_cpu.cpu.state.o_cnt[2] ),
    .A3(\u_cpu.cpu.mem_bytecnt[0] ),
    .ZN(_02338_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05856_ (.A1(\u_cpu.cpu.decode.op26 ),
    .A2(_01411_),
    .ZN(_02339_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _05857_ (.A1(_02337_),
    .A2(\u_cpu.cpu.state.o_cnt_r[3] ),
    .A3(_02338_),
    .A4(_02339_),
    .Z(_02340_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05858_ (.I(\u_cpu.cpu.genblk3.csr.mcause3_0[0] ),
    .ZN(_02341_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05859_ (.A1(_02311_),
    .A2(\u_cpu.cpu.genblk3.csr.mcause31 ),
    .B(_02338_),
    .ZN(_02342_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05860_ (.I(\u_cpu.cpu.decode.op21 ),
    .ZN(_02343_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _05861_ (.A1(_02343_),
    .A2(\u_cpu.cpu.decode.co_ebreak ),
    .A3(_01411_),
    .ZN(_02344_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05862_ (.A1(_02305_),
    .A2(_02344_),
    .ZN(_02345_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _05863_ (.A1(_02341_),
    .A2(_02338_),
    .B(_02342_),
    .C(_02345_),
    .ZN(_02346_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _05864_ (.A1(_02336_),
    .A2(_02324_),
    .B1(_02340_),
    .B2(\u_cpu.cpu.genblk3.csr.mstatus_mie ),
    .C(_02346_),
    .ZN(_02347_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _05865_ (.A1(_01409_),
    .A2(_02331_),
    .A3(_02334_),
    .B1(_02335_),
    .B2(_02347_),
    .ZN(_02348_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05866_ (.A1(_01393_),
    .A2(_02348_),
    .ZN(_02349_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05867_ (.A1(\u_arbiter.i_wb_cpu_ibus_adr[0] ),
    .A2(_01386_),
    .ZN(_02350_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05868_ (.A1(_02349_),
    .A2(_02350_),
    .ZN(\u_cpu.cpu.o_wdata1 ));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05869_ (.A1(_02309_),
    .A2(_02325_),
    .ZN(_02351_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05870_ (.A1(_02309_),
    .A2(_02325_),
    .B(_01369_),
    .ZN(_02352_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05871_ (.A1(\u_cpu.cpu.bne_or_bge ),
    .A2(_02351_),
    .B(_02352_),
    .ZN(_02353_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05872_ (.A1(_01370_),
    .A2(_02351_),
    .B(_02353_),
    .ZN(_02354_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05873_ (.I(\u_cpu.cpu.alu.cmp_r ),
    .ZN(_02355_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05874_ (.A1(\u_cpu.cpu.state.o_cnt_r[0] ),
    .A2(_02338_),
    .ZN(_02356_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _05875_ (.A1(_01369_),
    .A2(_02355_),
    .A3(_02356_),
    .ZN(_02357_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _05876_ (.A1(_02309_),
    .A2(\u_cpu.cpu.alu.add_cy_r ),
    .Z(_02358_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _05877_ (.A1(_02358_),
    .A2(_02308_),
    .A3(_02325_),
    .Z(_02359_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05878_ (.A1(_01410_),
    .A2(_02359_),
    .ZN(_02360_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05879_ (.I(\u_cpu.cpu.bufreg.lsb[0] ),
    .ZN(_02361_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _05880_ (.A1(_01384_),
    .A2(\u_cpu.cpu.state.init_done ),
    .A3(_01385_),
    .A4(_01375_),
    .ZN(_02362_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _05881_ (.A1(\u_cpu.cpu.branch_op ),
    .A2(_02313_),
    .Z(_02363_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _05882_ (.A1(_01369_),
    .A2(_01370_),
    .Z(_02364_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _05883_ (.A1(_01409_),
    .A2(_02363_),
    .A3(_02364_),
    .B(_01372_),
    .ZN(_02365_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _05884_ (.A1(_02305_),
    .A2(_02362_),
    .A3(_02365_),
    .ZN(_02366_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05885_ (.A1(_01373_),
    .A2(_01370_),
    .ZN(_02367_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05886_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[5] ),
    .A2(_01369_),
    .ZN(_02368_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05887_ (.A1(\u_cpu.cpu.state.stage_two_req ),
    .A2(_02368_),
    .ZN(_02369_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _05888_ (.A1(\u_cpu.cpu.state.init_done ),
    .A2(_02367_),
    .A3(_02369_),
    .ZN(_02370_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _05889_ (.A1(_02366_),
    .A2(_02370_),
    .Z(_02371_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05890_ (.I(_02371_),
    .Z(_02372_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05891_ (.A1(_02361_),
    .A2(_02372_),
    .ZN(_02373_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _05892_ (.A1(_01370_),
    .A2(_02357_),
    .B(_02360_),
    .C(_02373_),
    .ZN(_02374_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _05893_ (.A1(_02354_),
    .A2(_02374_),
    .B(_01373_),
    .C(_02363_),
    .ZN(_02375_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05894_ (.I(\u_cpu.cpu.state.o_cnt_r[1] ),
    .ZN(_02376_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05895_ (.A1(\u_cpu.cpu.state.o_cnt_r[2] ),
    .A2(\u_cpu.cpu.ctrl.i_iscomp ),
    .ZN(_02377_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05896_ (.A1(_02376_),
    .A2(\u_cpu.cpu.ctrl.i_iscomp ),
    .B(_02377_),
    .ZN(_02378_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _05897_ (.A1(_02338_),
    .A2(_02378_),
    .Z(_02379_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _05898_ (.A1(\u_arbiter.i_wb_cpu_ibus_adr[0] ),
    .A2(\u_cpu.cpu.ctrl.pc_plus_4_cy_r ),
    .Z(_02380_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _05899_ (.A1(_02379_),
    .A2(_02380_),
    .ZN(_02381_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05900_ (.A1(_01374_),
    .A2(_02313_),
    .ZN(_02382_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05901_ (.I(_02313_),
    .ZN(_02383_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05902_ (.I(\u_cpu.cpu.mem_if.signbit ),
    .ZN(_02384_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _05903_ (.A1(_02332_),
    .A2(\u_cpu.cpu.mem_bytecnt[1] ),
    .B1(\u_cpu.cpu.mem_bytecnt[0] ),
    .B2(_01409_),
    .ZN(_02385_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05904_ (.I0(\u_arbiter.i_wb_cpu_dbus_dat[0] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_dat[8] ),
    .I2(\u_arbiter.i_wb_cpu_dbus_dat[16] ),
    .I3(\u_arbiter.i_wb_cpu_dbus_dat[24] ),
    .S0(\u_cpu.cpu.bufreg.lsb[0] ),
    .S1(\u_cpu.cpu.bufreg.lsb[1] ),
    .Z(_02386_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05905_ (.A1(_02385_),
    .A2(_02386_),
    .ZN(_02387_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05906_ (.A1(_02384_),
    .A2(_02385_),
    .B(_02387_),
    .ZN(_00728_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05907_ (.A1(_01369_),
    .A2(_02387_),
    .ZN(_02388_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _05908_ (.A1(_01373_),
    .A2(_02383_),
    .A3(_00728_),
    .A4(_02388_),
    .ZN(_02389_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _05909_ (.A1(_02381_),
    .A2(_02382_),
    .B(_02347_),
    .C(_02389_),
    .ZN(_02390_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05910_ (.A1(_01372_),
    .A2(_02313_),
    .ZN(_02391_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _05911_ (.A1(\u_cpu.cpu.immdec.imm31 ),
    .A2(_02317_),
    .Z(_02392_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _05912_ (.A1(_02311_),
    .A2(_02315_),
    .A3(_02316_),
    .ZN(_02393_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05913_ (.A1(_02311_),
    .A2(_02392_),
    .B(_02393_),
    .ZN(_02394_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _05914_ (.A1(\u_cpu.cpu.state.o_cnt[2] ),
    .A2(\u_cpu.cpu.mem_bytecnt[0] ),
    .Z(_02395_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05915_ (.A1(_01374_),
    .A2(_02391_),
    .ZN(_02396_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05916_ (.A1(\u_cpu.cpu.mem_bytecnt[1] ),
    .A2(_02395_),
    .B(_02396_),
    .ZN(_02397_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05917_ (.A1(_02394_),
    .A2(_02397_),
    .ZN(_02398_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _05918_ (.A1(_02361_),
    .A2(_02396_),
    .A3(_02372_),
    .ZN(_02399_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05919_ (.A1(\u_cpu.cpu.decode.opcode[1] ),
    .A2(_02313_),
    .B(_02314_),
    .ZN(_02400_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _05920_ (.A1(_01374_),
    .A2(_02306_),
    .B1(_01381_),
    .B2(_01378_),
    .C(_02400_),
    .ZN(_02401_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05921_ (.A1(\u_arbiter.i_wb_cpu_ibus_adr[0] ),
    .A2(_02401_),
    .ZN(_02402_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _05922_ (.A1(\u_cpu.cpu.ctrl.pc_plus_offset_cy_r ),
    .A2(_02402_),
    .ZN(_02403_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05923_ (.A1(_02398_),
    .A2(_02399_),
    .B(_02403_),
    .ZN(_02404_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _05924_ (.A1(_02403_),
    .A2(_02398_),
    .A3(_02399_),
    .Z(_02405_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _05925_ (.A1(_02404_),
    .A2(_02356_),
    .A3(_02405_),
    .ZN(_02406_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _05926_ (.A1(_01374_),
    .A2(_02391_),
    .A3(_02406_),
    .ZN(_02407_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _05927_ (.A1(_02375_),
    .A2(_02390_),
    .A3(_02407_),
    .ZN(_02408_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05928_ (.A1(_01374_),
    .A2(_02406_),
    .ZN(_02409_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _05929_ (.A1(_01374_),
    .A2(_02373_),
    .B(_02409_),
    .C(_01386_),
    .ZN(_02410_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05930_ (.A1(_01386_),
    .A2(_02408_),
    .B(_02410_),
    .ZN(_02411_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05931_ (.I(_02411_),
    .Z(\u_cpu.cpu.o_wdata0 ));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05932_ (.A1(_02321_),
    .A2(\u_cpu.rf_ram.rdata[1] ),
    .ZN(_02412_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05933_ (.A1(_02320_),
    .A2(\u_cpu.rf_ram_if.rdata1[1] ),
    .ZN(_02413_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05934_ (.A1(_02320_),
    .A2(_02412_),
    .B(_02413_),
    .ZN(_00015_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05935_ (.A1(_02321_),
    .A2(\u_cpu.rf_ram.rdata[2] ),
    .ZN(_02414_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05936_ (.A1(_02320_),
    .A2(\u_cpu.rf_ram_if.rdata1[2] ),
    .ZN(_02415_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05937_ (.A1(_02320_),
    .A2(_02414_),
    .B(_02415_),
    .ZN(_00016_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05938_ (.A1(_02321_),
    .A2(\u_cpu.rf_ram.rdata[3] ),
    .ZN(_02416_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05939_ (.A1(_02320_),
    .A2(\u_cpu.rf_ram_if.rdata1[3] ),
    .ZN(_02417_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05940_ (.A1(_02320_),
    .A2(_02416_),
    .B(_02417_),
    .ZN(_00017_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05941_ (.A1(_02321_),
    .A2(\u_cpu.rf_ram.rdata[4] ),
    .ZN(_02418_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05942_ (.A1(_02320_),
    .A2(\u_cpu.rf_ram_if.rdata1[4] ),
    .ZN(_02419_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05943_ (.A1(_02320_),
    .A2(_02418_),
    .B(_02419_),
    .ZN(_00018_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05944_ (.A1(_02321_),
    .A2(\u_cpu.rf_ram.rdata[5] ),
    .ZN(_02420_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05945_ (.A1(_02320_),
    .A2(\u_cpu.rf_ram_if.rdata1[5] ),
    .ZN(_02421_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05946_ (.A1(_02320_),
    .A2(_02420_),
    .B(_02421_),
    .ZN(_00019_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05947_ (.A1(_02321_),
    .A2(\u_cpu.rf_ram.rdata[6] ),
    .ZN(_02422_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05948_ (.A1(_02320_),
    .A2(\u_cpu.rf_ram_if.rdata1[6] ),
    .ZN(_02423_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05949_ (.A1(_02320_),
    .A2(_02422_),
    .B(_02423_),
    .ZN(_00020_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05950_ (.A1(\u_cpu.rf_ram_if.rdata0[1] ),
    .A2(_01403_),
    .ZN(_02424_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05951_ (.A1(_01403_),
    .A2(_02322_),
    .B(_02424_),
    .ZN(_00008_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05952_ (.A1(\u_cpu.rf_ram_if.rdata0[2] ),
    .A2(_01403_),
    .ZN(_02425_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05953_ (.A1(_01403_),
    .A2(_02412_),
    .B(_02425_),
    .ZN(_00009_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05954_ (.A1(\u_cpu.rf_ram_if.rdata0[3] ),
    .A2(_01403_),
    .ZN(_02426_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05955_ (.A1(_01403_),
    .A2(_02414_),
    .B(_02426_),
    .ZN(_00010_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05956_ (.A1(\u_cpu.rf_ram_if.rdata0[4] ),
    .A2(_01403_),
    .ZN(_02427_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05957_ (.A1(_01403_),
    .A2(_02416_),
    .B(_02427_),
    .ZN(_00011_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05958_ (.A1(\u_cpu.rf_ram_if.rdata0[5] ),
    .A2(_01403_),
    .ZN(_02428_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05959_ (.A1(_01403_),
    .A2(_02418_),
    .B(_02428_),
    .ZN(_00012_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05960_ (.A1(\u_cpu.rf_ram_if.rdata0[6] ),
    .A2(_01403_),
    .ZN(_02429_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05961_ (.A1(_01403_),
    .A2(_02420_),
    .B(_02429_),
    .ZN(_00013_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05962_ (.A1(\u_cpu.rf_ram_if.rdata0[7] ),
    .A2(_01403_),
    .ZN(_02430_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05963_ (.A1(_01403_),
    .A2(_02422_),
    .B(_02430_),
    .ZN(_00014_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05964_ (.I(\u_cpu.cpu.bufreg.lsb[1] ),
    .ZN(_02431_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _05965_ (.A1(_02332_),
    .A2(_02431_),
    .B1(_01409_),
    .B2(_02361_),
    .ZN(_02432_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _05966_ (.A1(\u_cpu.cpu.state.o_cnt_r[0] ),
    .A2(\u_cpu.cpu.state.o_cnt_r[1] ),
    .A3(\u_cpu.cpu.state.o_cnt_r[2] ),
    .A4(\u_cpu.cpu.state.o_cnt_r[3] ),
    .ZN(_02433_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05967_ (.A1(_01372_),
    .A2(_01374_),
    .ZN(_02434_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _05968_ (.A1(\u_cpu.cpu.state.init_done ),
    .A2(_02433_),
    .A3(_02434_),
    .ZN(_02435_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05969_ (.A1(_02432_),
    .A2(_02435_),
    .B(_01445_),
    .ZN(\u_arbiter.o_wb_cpu_cyc ));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05970_ (.I(_02306_),
    .ZN(_02436_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05971_ (.A1(_02436_),
    .A2(_01431_),
    .ZN(\u_arbiter.o_wb_cpu_we ));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05972_ (.A1(_01374_),
    .A2(\u_cpu.cpu.decode.opcode[1] ),
    .ZN(_02437_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05973_ (.A1(_01374_),
    .A2(_02383_),
    .ZN(_02438_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _05974_ (.A1(_02309_),
    .A2(\u_cpu.cpu.bufreg.c_r ),
    .A3(_02437_),
    .A4(_02438_),
    .ZN(_02439_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _05975_ (.A1(\u_cpu.cpu.decode.opcode[1] ),
    .A2(_02313_),
    .Z(_02440_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _05976_ (.A1(_01375_),
    .A2(_02356_),
    .A3(_02440_),
    .ZN(_02441_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _05977_ (.A1(_02309_),
    .A2(_02437_),
    .A3(_02438_),
    .ZN(_02442_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _05978_ (.A1(\u_cpu.cpu.bufreg.c_r ),
    .A2(_02442_),
    .Z(_02443_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _05979_ (.A1(_01372_),
    .A2(_02394_),
    .A3(_02441_),
    .A4(_02443_),
    .Z(_02444_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05980_ (.I(_02372_),
    .Z(_02445_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05981_ (.A1(_02439_),
    .A2(_02444_),
    .B(_02445_),
    .ZN(_00022_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _05982_ (.A1(\u_arbiter.i_wb_cpu_ibus_adr[0] ),
    .A2(\u_cpu.cpu.ctrl.pc_plus_offset_cy_r ),
    .A3(_02401_),
    .ZN(_02446_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05983_ (.A1(\u_cpu.cpu.genblk3.csr.o_new_irq ),
    .A2(\u_cpu.cpu.state.init_done ),
    .ZN(_02447_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05984_ (.A1(_02447_),
    .A2(_02365_),
    .ZN(_02448_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05985_ (.A1(_02305_),
    .A2(_02448_),
    .ZN(_02449_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05986_ (.A1(_02446_),
    .A2(_02404_),
    .B(_02449_),
    .ZN(_00024_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05987_ (.A1(\u_arbiter.i_wb_cpu_ibus_adr[0] ),
    .A2(\u_cpu.cpu.ctrl.pc_plus_4_cy_r ),
    .ZN(_02450_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05988_ (.A1(_02379_),
    .A2(_02380_),
    .ZN(_02451_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05989_ (.A1(_02450_),
    .A2(_02451_),
    .B(_02449_),
    .ZN(_00023_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05990_ (.A1(_01387_),
    .A2(_02433_),
    .ZN(\u_cpu.cpu.o_wen1 ));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _05991_ (.A1(\u_cpu.cpu.immdec.imm11_7[1] ),
    .A2(\u_cpu.cpu.immdec.imm11_7[2] ),
    .A3(\u_cpu.cpu.immdec.imm11_7[3] ),
    .A4(\u_cpu.cpu.immdec.imm11_7[0] ),
    .Z(_02452_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _05992_ (.A1(_02306_),
    .A2(_02313_),
    .B(_02382_),
    .C(_01373_),
    .ZN(_02453_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _05993_ (.A1(\u_cpu.cpu.immdec.imm11_7[4] ),
    .A2(_02452_),
    .B(_02453_),
    .C(_02448_),
    .ZN(_02454_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05994_ (.A1(_01393_),
    .A2(_02454_),
    .B(_02433_),
    .ZN(\u_cpu.cpu.o_wen0 ));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05995_ (.A1(\u_cpu.cpu.bufreg.lsb[0] ),
    .A2(\u_cpu.cpu.bne_or_bge ),
    .ZN(_02455_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05996_ (.A1(\u_cpu.cpu.bufreg.lsb[1] ),
    .A2(_02455_),
    .B(_02332_),
    .ZN(\u_arbiter.i_wb_cpu_dbus_sel[1] ));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05997_ (.A1(\u_cpu.cpu.bufreg.lsb[0] ),
    .A2(_02431_),
    .B(_02332_),
    .ZN(\u_arbiter.i_wb_cpu_dbus_sel[2] ));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05998_ (.A1(_02431_),
    .A2(_02455_),
    .B(_02332_),
    .ZN(\u_arbiter.i_wb_cpu_dbus_sel[3] ));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05999_ (.A1(_01386_),
    .A2(_01394_),
    .B(\u_cpu.rf_ram_if.genblk1.wtrig0_r ),
    .ZN(_02456_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06000_ (.A1(\u_cpu.rf_ram_if.genblk1.wtrig0_r ),
    .A2(_01386_),
    .ZN(_02457_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06001_ (.A1(_02312_),
    .A2(_02457_),
    .ZN(_02458_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06002_ (.A1(_02456_),
    .A2(_02458_),
    .ZN(_02459_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _06003_ (.I(\u_cpu.rf_ram_if.genblk1.wtrig0_r ),
    .ZN(_02460_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06004_ (.A1(\u_cpu.cpu.immdec.imm11_7[1] ),
    .A2(_02460_),
    .ZN(_02461_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06005_ (.A1(_02460_),
    .A2(_01412_),
    .B(_02461_),
    .ZN(_02462_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06006_ (.A1(_01386_),
    .A2(_02462_),
    .ZN(_02463_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06007_ (.A1(_02459_),
    .A2(_02463_),
    .ZN(_02464_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06008_ (.A1(\u_cpu.rf_ram_if.rcnt[1] ),
    .A2(\u_cpu.rf_ram_if.rcnt[0] ),
    .B(\u_cpu.rf_ram_if.rcnt[2] ),
    .ZN(_02465_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06009_ (.A1(_01543_),
    .A2(_02465_),
    .Z(_02466_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06010_ (.I(_02466_),
    .ZN(_02467_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06011_ (.A1(_01591_),
    .A2(_02467_),
    .ZN(_02468_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06012_ (.A1(_02464_),
    .A2(_02468_),
    .ZN(_02469_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06013_ (.A1(\u_cpu.cpu.immdec.imm11_7[2] ),
    .A2(_02457_),
    .ZN(_02470_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06014_ (.A1(\u_cpu.rf_ram_if.genblk1.wtrig0_r ),
    .A2(\u_cpu.rf_ram_if.wen1_r ),
    .B1(\u_cpu.rf_ram_if.rtrig0 ),
    .B2(\u_cpu.rf_ram_if.wen0_r ),
    .ZN(_02471_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06015_ (.I(_02471_),
    .ZN(_02472_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06016_ (.A1(\u_cpu.cpu.immdec.imm11_7[4] ),
    .A2(_02457_),
    .A3(_02472_),
    .ZN(_02473_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _06017_ (.A1(\u_cpu.cpu.immdec.imm11_7[3] ),
    .A2(_02470_),
    .A3(_02473_),
    .ZN(_02474_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06018_ (.I(_02474_),
    .Z(_02475_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06019_ (.A1(_02469_),
    .A2(_02475_),
    .ZN(_02476_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06020_ (.I(_02476_),
    .Z(_02477_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06021_ (.I(\u_cpu.rf_ram_if.genblk1.wtrig0_r ),
    .Z(_02478_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06022_ (.A1(\u_cpu.rf_ram_if.wdata1_r[0] ),
    .A2(_02478_),
    .Z(_02479_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06023_ (.A1(\u_cpu.rf_ram_if.wdata0_r[0] ),
    .A2(_02460_),
    .B(_02479_),
    .ZN(_02480_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06024_ (.I(_02480_),
    .Z(_02481_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06025_ (.I(_02481_),
    .Z(_02482_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06026_ (.A1(\u_cpu.rf_ram.memory[82][0] ),
    .A2(_02477_),
    .ZN(_02483_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06027_ (.A1(_02477_),
    .A2(_02482_),
    .B(_02483_),
    .ZN(_00026_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06028_ (.A1(_02478_),
    .A2(\u_cpu.rf_ram_if.wdata1_r[1] ),
    .Z(_02484_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06029_ (.A1(_02460_),
    .A2(\u_cpu.rf_ram_if.wdata0_r[1] ),
    .B(_02484_),
    .ZN(_02485_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06030_ (.I(_02485_),
    .Z(_02486_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06031_ (.I(_02486_),
    .Z(_02487_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06032_ (.A1(\u_cpu.rf_ram.memory[82][1] ),
    .A2(_02477_),
    .ZN(_02488_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06033_ (.A1(_02477_),
    .A2(_02487_),
    .B(_02488_),
    .ZN(_00027_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06034_ (.A1(_02478_),
    .A2(\u_cpu.rf_ram_if.wdata1_r[2] ),
    .Z(_02489_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06035_ (.A1(_02460_),
    .A2(\u_cpu.rf_ram_if.wdata0_r[2] ),
    .B(_02489_),
    .ZN(_02490_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06036_ (.I(_02490_),
    .Z(_02491_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06037_ (.I(_02491_),
    .Z(_02492_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06038_ (.A1(\u_cpu.rf_ram.memory[82][2] ),
    .A2(_02477_),
    .ZN(_02493_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06039_ (.A1(_02477_),
    .A2(_02492_),
    .B(_02493_),
    .ZN(_00028_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06040_ (.A1(_02478_),
    .A2(\u_cpu.rf_ram_if.wdata1_r[3] ),
    .Z(_02494_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06041_ (.A1(_02460_),
    .A2(\u_cpu.rf_ram_if.wdata0_r[3] ),
    .B(_02494_),
    .ZN(_02495_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06042_ (.I(_02495_),
    .Z(_02496_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06043_ (.I(_02496_),
    .Z(_02497_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06044_ (.A1(\u_cpu.rf_ram.memory[82][3] ),
    .A2(_02477_),
    .ZN(_02498_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06045_ (.A1(_02477_),
    .A2(_02497_),
    .B(_02498_),
    .ZN(_00029_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06046_ (.A1(_02478_),
    .A2(\u_cpu.rf_ram_if.wdata1_r[4] ),
    .Z(_02499_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06047_ (.A1(_02460_),
    .A2(\u_cpu.rf_ram_if.wdata0_r[4] ),
    .B(_02499_),
    .ZN(_02500_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06048_ (.I(_02500_),
    .Z(_02501_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06049_ (.I(_02501_),
    .Z(_02502_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06050_ (.A1(\u_cpu.rf_ram.memory[82][4] ),
    .A2(_02477_),
    .ZN(_02503_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06051_ (.A1(_02477_),
    .A2(_02502_),
    .B(_02503_),
    .ZN(_00030_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06052_ (.A1(_02478_),
    .A2(\u_cpu.rf_ram_if.wdata1_r[5] ),
    .Z(_02504_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06053_ (.A1(_02460_),
    .A2(\u_cpu.rf_ram_if.wdata0_r[5] ),
    .B(_02504_),
    .ZN(_02505_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06054_ (.I(_02505_),
    .Z(_02506_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06055_ (.I(_02506_),
    .Z(_02507_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06056_ (.A1(\u_cpu.rf_ram.memory[82][5] ),
    .A2(_02477_),
    .ZN(_02508_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06057_ (.A1(_02477_),
    .A2(_02507_),
    .B(_02508_),
    .ZN(_00031_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06058_ (.A1(_02478_),
    .A2(\u_cpu.rf_ram_if.wdata1_r[6] ),
    .Z(_02509_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06059_ (.A1(_02460_),
    .A2(\u_cpu.rf_ram_if.wdata0_r[6] ),
    .B(_02509_),
    .ZN(_02510_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06060_ (.I(_02510_),
    .Z(_02511_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06061_ (.I(_02511_),
    .Z(_02512_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06062_ (.A1(\u_cpu.rf_ram.memory[82][6] ),
    .A2(_02477_),
    .ZN(_02513_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06063_ (.A1(_02477_),
    .A2(_02512_),
    .B(_02513_),
    .ZN(_00032_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06064_ (.A1(_02478_),
    .A2(\u_cpu.rf_ram_if.wdata1_r[7] ),
    .Z(_02514_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06065_ (.A1(_02460_),
    .A2(\u_cpu.cpu.o_wdata0 ),
    .B(_02514_),
    .ZN(_02515_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06066_ (.I(_02515_),
    .Z(_02516_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06067_ (.I(_02516_),
    .Z(_02517_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06068_ (.A1(\u_cpu.rf_ram.memory[82][7] ),
    .A2(_02477_),
    .ZN(_02518_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06069_ (.A1(_02477_),
    .A2(_02517_),
    .B(_02518_),
    .ZN(_00033_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _06070_ (.A1(\u_cpu.rf_ram_if.rcnt[1] ),
    .A2(\u_cpu.rf_ram_if.rcnt[0] ),
    .B(_01543_),
    .C(\u_cpu.rf_ram_if.rcnt[2] ),
    .ZN(_02519_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06071_ (.A1(_01547_),
    .A2(_02519_),
    .Z(_02520_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _06072_ (.A1(_02467_),
    .A2(_02520_),
    .Z(_02521_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06073_ (.A1(_02456_),
    .A2(_02458_),
    .Z(_02522_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06074_ (.A1(_02522_),
    .A2(_02463_),
    .ZN(_02523_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06075_ (.A1(_02521_),
    .A2(_02523_),
    .ZN(_02524_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06076_ (.I(\u_cpu.cpu.immdec.imm11_7[4] ),
    .ZN(_02525_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06077_ (.A1(_02525_),
    .A2(_02472_),
    .ZN(_02526_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _06078_ (.A1(\u_cpu.cpu.immdec.imm11_7[3] ),
    .A2(_02470_),
    .A3(_02526_),
    .ZN(_02527_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06079_ (.I(_02527_),
    .Z(_02528_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06080_ (.A1(_02524_),
    .A2(_02528_),
    .ZN(_02529_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06081_ (.I(_02529_),
    .Z(_02530_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06082_ (.A1(\u_cpu.rf_ram.memory[21][0] ),
    .A2(_02530_),
    .ZN(_02531_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06083_ (.A1(_02482_),
    .A2(_02530_),
    .B(_02531_),
    .ZN(_00034_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06084_ (.A1(\u_cpu.rf_ram.memory[21][1] ),
    .A2(_02530_),
    .ZN(_02532_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06085_ (.A1(_02487_),
    .A2(_02530_),
    .B(_02532_),
    .ZN(_00035_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06086_ (.A1(\u_cpu.rf_ram.memory[21][2] ),
    .A2(_02530_),
    .ZN(_02533_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06087_ (.A1(_02492_),
    .A2(_02530_),
    .B(_02533_),
    .ZN(_00036_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06088_ (.A1(\u_cpu.rf_ram.memory[21][3] ),
    .A2(_02530_),
    .ZN(_02534_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06089_ (.A1(_02497_),
    .A2(_02530_),
    .B(_02534_),
    .ZN(_00037_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06090_ (.A1(\u_cpu.rf_ram.memory[21][4] ),
    .A2(_02530_),
    .ZN(_02535_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06091_ (.A1(_02502_),
    .A2(_02530_),
    .B(_02535_),
    .ZN(_00038_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06092_ (.A1(\u_cpu.rf_ram.memory[21][5] ),
    .A2(_02530_),
    .ZN(_02536_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06093_ (.A1(_02507_),
    .A2(_02530_),
    .B(_02536_),
    .ZN(_00039_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06094_ (.A1(\u_cpu.rf_ram.memory[21][6] ),
    .A2(_02530_),
    .ZN(_02537_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06095_ (.A1(_02512_),
    .A2(_02530_),
    .B(_02537_),
    .ZN(_00040_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06096_ (.A1(\u_cpu.rf_ram.memory[21][7] ),
    .A2(_02530_),
    .ZN(_02538_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06097_ (.A1(_02517_),
    .A2(_02530_),
    .B(_02538_),
    .ZN(_00041_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06098_ (.A1(_02464_),
    .A2(_02521_),
    .ZN(_02539_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06099_ (.A1(_02475_),
    .A2(_02539_),
    .ZN(_02540_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06100_ (.I(_02540_),
    .Z(_02541_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06101_ (.A1(\u_cpu.rf_ram.memory[81][0] ),
    .A2(_02541_),
    .ZN(_02542_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06102_ (.A1(_02482_),
    .A2(_02541_),
    .B(_02542_),
    .ZN(_00042_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06103_ (.A1(\u_cpu.rf_ram.memory[81][1] ),
    .A2(_02541_),
    .ZN(_02543_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06104_ (.A1(_02487_),
    .A2(_02541_),
    .B(_02543_),
    .ZN(_00043_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06105_ (.A1(\u_cpu.rf_ram.memory[81][2] ),
    .A2(_02541_),
    .ZN(_02544_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06106_ (.A1(_02492_),
    .A2(_02541_),
    .B(_02544_),
    .ZN(_00044_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06107_ (.A1(\u_cpu.rf_ram.memory[81][3] ),
    .A2(_02541_),
    .ZN(_02545_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06108_ (.A1(_02497_),
    .A2(_02541_),
    .B(_02545_),
    .ZN(_00045_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06109_ (.A1(\u_cpu.rf_ram.memory[81][4] ),
    .A2(_02541_),
    .ZN(_02546_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06110_ (.A1(_02502_),
    .A2(_02541_),
    .B(_02546_),
    .ZN(_00046_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06111_ (.A1(\u_cpu.rf_ram.memory[81][5] ),
    .A2(_02541_),
    .ZN(_02547_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06112_ (.A1(_02507_),
    .A2(_02541_),
    .B(_02547_),
    .ZN(_00047_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06113_ (.A1(\u_cpu.rf_ram.memory[81][6] ),
    .A2(_02541_),
    .ZN(_02548_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06114_ (.A1(_02512_),
    .A2(_02541_),
    .B(_02548_),
    .ZN(_00048_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06115_ (.A1(\u_cpu.rf_ram.memory[81][7] ),
    .A2(_02541_),
    .ZN(_02549_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06116_ (.A1(_02517_),
    .A2(_02541_),
    .B(_02549_),
    .ZN(_00049_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06117_ (.A1(_02469_),
    .A2(_02528_),
    .ZN(_02550_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06118_ (.I(_02550_),
    .Z(_02551_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06119_ (.A1(\u_cpu.rf_ram.memory[18][0] ),
    .A2(_02551_),
    .ZN(_02552_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06120_ (.A1(_02482_),
    .A2(_02551_),
    .B(_02552_),
    .ZN(_00050_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06121_ (.A1(\u_cpu.rf_ram.memory[18][1] ),
    .A2(_02551_),
    .ZN(_02553_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06122_ (.A1(_02487_),
    .A2(_02551_),
    .B(_02553_),
    .ZN(_00051_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06123_ (.A1(\u_cpu.rf_ram.memory[18][2] ),
    .A2(_02551_),
    .ZN(_02554_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06124_ (.A1(_02492_),
    .A2(_02551_),
    .B(_02554_),
    .ZN(_00052_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06125_ (.A1(\u_cpu.rf_ram.memory[18][3] ),
    .A2(_02551_),
    .ZN(_02555_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06126_ (.A1(_02497_),
    .A2(_02551_),
    .B(_02555_),
    .ZN(_00053_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06127_ (.A1(\u_cpu.rf_ram.memory[18][4] ),
    .A2(_02551_),
    .ZN(_02556_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06128_ (.A1(_02502_),
    .A2(_02551_),
    .B(_02556_),
    .ZN(_00054_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06129_ (.A1(\u_cpu.rf_ram.memory[18][5] ),
    .A2(_02551_),
    .ZN(_02557_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06130_ (.A1(_02507_),
    .A2(_02551_),
    .B(_02557_),
    .ZN(_00055_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06131_ (.A1(\u_cpu.rf_ram.memory[18][6] ),
    .A2(_02551_),
    .ZN(_02558_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06132_ (.A1(_02512_),
    .A2(_02551_),
    .B(_02558_),
    .ZN(_00056_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06133_ (.A1(\u_cpu.rf_ram.memory[18][7] ),
    .A2(_02551_),
    .ZN(_02559_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06134_ (.A1(_02517_),
    .A2(_02551_),
    .B(_02559_),
    .ZN(_00057_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _06135_ (.A1(_01668_),
    .A2(_02466_),
    .Z(_02560_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06136_ (.A1(_02523_),
    .A2(_02560_),
    .ZN(_02561_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06137_ (.A1(_02528_),
    .A2(_02561_),
    .ZN(_02562_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06138_ (.I(_02562_),
    .Z(_02563_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06139_ (.A1(\u_cpu.rf_ram.memory[20][0] ),
    .A2(_02563_),
    .ZN(_02564_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06140_ (.A1(_02482_),
    .A2(_02563_),
    .B(_02564_),
    .ZN(_00058_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06141_ (.A1(\u_cpu.rf_ram.memory[20][1] ),
    .A2(_02563_),
    .ZN(_02565_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06142_ (.A1(_02487_),
    .A2(_02563_),
    .B(_02565_),
    .ZN(_00059_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06143_ (.A1(\u_cpu.rf_ram.memory[20][2] ),
    .A2(_02563_),
    .ZN(_02566_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06144_ (.A1(_02492_),
    .A2(_02563_),
    .B(_02566_),
    .ZN(_00060_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06145_ (.A1(\u_cpu.rf_ram.memory[20][3] ),
    .A2(_02563_),
    .ZN(_02567_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06146_ (.A1(_02497_),
    .A2(_02563_),
    .B(_02567_),
    .ZN(_00061_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06147_ (.A1(\u_cpu.rf_ram.memory[20][4] ),
    .A2(_02563_),
    .ZN(_02568_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06148_ (.A1(_02502_),
    .A2(_02563_),
    .B(_02568_),
    .ZN(_00062_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06149_ (.A1(\u_cpu.rf_ram.memory[20][5] ),
    .A2(_02563_),
    .ZN(_02569_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06150_ (.A1(_02507_),
    .A2(_02563_),
    .B(_02569_),
    .ZN(_00063_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06151_ (.A1(\u_cpu.rf_ram.memory[20][6] ),
    .A2(_02563_),
    .ZN(_02570_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06152_ (.A1(_02512_),
    .A2(_02563_),
    .B(_02570_),
    .ZN(_00064_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06153_ (.A1(\u_cpu.rf_ram.memory[20][7] ),
    .A2(_02563_),
    .ZN(_02571_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06154_ (.A1(_02517_),
    .A2(_02563_),
    .B(_02571_),
    .ZN(_00065_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06155_ (.I0(\u_cpu.rf_ram_if.wdata0_r[0] ),
    .I1(\u_cpu.rf_ram_if.wdata1_r[0] ),
    .S(_02478_),
    .Z(_02572_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06156_ (.I(_02572_),
    .Z(_02573_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06157_ (.A1(\u_cpu.cpu.immdec.imm11_7[3] ),
    .A2(_02457_),
    .ZN(_02574_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06158_ (.A1(_02470_),
    .A2(_02574_),
    .ZN(_02575_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _06159_ (.A1(_02478_),
    .A2(_01386_),
    .A3(_02526_),
    .A4(_02575_),
    .ZN(_02576_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06160_ (.I(_02576_),
    .Z(_02577_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06161_ (.A1(_02539_),
    .A2(_02577_),
    .ZN(_02578_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06162_ (.I0(_02573_),
    .I1(\u_cpu.rf_ram.memory[1][0] ),
    .S(_02578_),
    .Z(_02579_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06163_ (.I(_02579_),
    .Z(_00066_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06164_ (.I0(\u_cpu.rf_ram_if.wdata0_r[1] ),
    .I1(\u_cpu.rf_ram_if.wdata1_r[1] ),
    .S(_02478_),
    .Z(_02580_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06165_ (.I(_02580_),
    .Z(_02581_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06166_ (.I0(_02581_),
    .I1(\u_cpu.rf_ram.memory[1][1] ),
    .S(_02578_),
    .Z(_02582_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06167_ (.I(_02582_),
    .Z(_00067_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06168_ (.I0(\u_cpu.rf_ram_if.wdata0_r[2] ),
    .I1(\u_cpu.rf_ram_if.wdata1_r[2] ),
    .S(_02478_),
    .Z(_02583_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06169_ (.I(_02583_),
    .Z(_02584_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06170_ (.I0(_02584_),
    .I1(\u_cpu.rf_ram.memory[1][2] ),
    .S(_02578_),
    .Z(_02585_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06171_ (.I(_02585_),
    .Z(_00068_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06172_ (.I0(\u_cpu.rf_ram_if.wdata0_r[3] ),
    .I1(\u_cpu.rf_ram_if.wdata1_r[3] ),
    .S(_02478_),
    .Z(_02586_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06173_ (.I(_02586_),
    .Z(_02587_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06174_ (.I0(_02587_),
    .I1(\u_cpu.rf_ram.memory[1][3] ),
    .S(_02578_),
    .Z(_02588_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06175_ (.I(_02588_),
    .Z(_00069_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06176_ (.I0(\u_cpu.rf_ram_if.wdata0_r[4] ),
    .I1(\u_cpu.rf_ram_if.wdata1_r[4] ),
    .S(_02478_),
    .Z(_02589_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06177_ (.I(_02589_),
    .Z(_02590_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06178_ (.I0(_02590_),
    .I1(\u_cpu.rf_ram.memory[1][4] ),
    .S(_02578_),
    .Z(_02591_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06179_ (.I(_02591_),
    .Z(_00070_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06180_ (.I0(\u_cpu.rf_ram_if.wdata0_r[5] ),
    .I1(\u_cpu.rf_ram_if.wdata1_r[5] ),
    .S(_02478_),
    .Z(_02592_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06181_ (.I(_02592_),
    .Z(_02593_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06182_ (.I0(_02593_),
    .I1(\u_cpu.rf_ram.memory[1][5] ),
    .S(_02578_),
    .Z(_02594_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06183_ (.I(_02594_),
    .Z(_00071_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06184_ (.I0(\u_cpu.rf_ram_if.wdata0_r[6] ),
    .I1(\u_cpu.rf_ram_if.wdata1_r[6] ),
    .S(_02478_),
    .Z(_02595_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06185_ (.I(_02595_),
    .Z(_02596_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06186_ (.I0(_02596_),
    .I1(\u_cpu.rf_ram.memory[1][6] ),
    .S(_02578_),
    .Z(_02597_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06187_ (.I(_02597_),
    .Z(_00072_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06188_ (.I0(\u_cpu.rf_ram_if.wdata1_r[7] ),
    .I1(\u_cpu.cpu.o_wdata0 ),
    .S(_02460_),
    .Z(_02598_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06189_ (.I(_02598_),
    .Z(_02599_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06190_ (.I0(_02599_),
    .I1(\u_cpu.rf_ram.memory[1][7] ),
    .S(_02578_),
    .Z(_02600_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06191_ (.I(_02600_),
    .Z(_00073_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06192_ (.A1(_02466_),
    .A2(_02520_),
    .ZN(_02601_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06193_ (.A1(_02523_),
    .A2(_02601_),
    .ZN(_02602_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06194_ (.A1(_02577_),
    .A2(_02602_),
    .ZN(_02603_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06195_ (.I0(_02573_),
    .I1(\u_cpu.rf_ram.memory[7][0] ),
    .S(_02603_),
    .Z(_02604_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06196_ (.I(_02604_),
    .Z(_00074_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06197_ (.I0(_02581_),
    .I1(\u_cpu.rf_ram.memory[7][1] ),
    .S(_02603_),
    .Z(_02605_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06198_ (.I(_02605_),
    .Z(_00075_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06199_ (.I0(_02584_),
    .I1(\u_cpu.rf_ram.memory[7][2] ),
    .S(_02603_),
    .Z(_02606_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06200_ (.I(_02606_),
    .Z(_00076_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06201_ (.I0(_02587_),
    .I1(\u_cpu.rf_ram.memory[7][3] ),
    .S(_02603_),
    .Z(_02607_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06202_ (.I(_02607_),
    .Z(_00077_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06203_ (.I0(_02590_),
    .I1(\u_cpu.rf_ram.memory[7][4] ),
    .S(_02603_),
    .Z(_02608_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06204_ (.I(_02608_),
    .Z(_00078_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06205_ (.I0(_02593_),
    .I1(\u_cpu.rf_ram.memory[7][5] ),
    .S(_02603_),
    .Z(_02609_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06206_ (.I(_02609_),
    .Z(_00079_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06207_ (.I0(_02596_),
    .I1(\u_cpu.rf_ram.memory[7][6] ),
    .S(_02603_),
    .Z(_02610_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06208_ (.I(_02610_),
    .Z(_00080_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06209_ (.I0(_02599_),
    .I1(\u_cpu.rf_ram.memory[7][7] ),
    .S(_02603_),
    .Z(_02611_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06210_ (.I(_02611_),
    .Z(_00081_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06211_ (.A1(_02464_),
    .A2(_02560_),
    .ZN(_02612_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06212_ (.A1(_02475_),
    .A2(_02612_),
    .ZN(_02613_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06213_ (.I(_02613_),
    .Z(_02614_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06214_ (.A1(\u_cpu.rf_ram.memory[80][0] ),
    .A2(_02614_),
    .ZN(_02615_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06215_ (.A1(_02482_),
    .A2(_02614_),
    .B(_02615_),
    .ZN(_00082_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06216_ (.A1(\u_cpu.rf_ram.memory[80][1] ),
    .A2(_02614_),
    .ZN(_02616_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06217_ (.A1(_02487_),
    .A2(_02614_),
    .B(_02616_),
    .ZN(_00083_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06218_ (.A1(\u_cpu.rf_ram.memory[80][2] ),
    .A2(_02614_),
    .ZN(_02617_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06219_ (.A1(_02492_),
    .A2(_02614_),
    .B(_02617_),
    .ZN(_00084_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06220_ (.A1(\u_cpu.rf_ram.memory[80][3] ),
    .A2(_02614_),
    .ZN(_02618_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06221_ (.A1(_02497_),
    .A2(_02614_),
    .B(_02618_),
    .ZN(_00085_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06222_ (.A1(\u_cpu.rf_ram.memory[80][4] ),
    .A2(_02614_),
    .ZN(_02619_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06223_ (.A1(_02502_),
    .A2(_02614_),
    .B(_02619_),
    .ZN(_00086_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06224_ (.A1(\u_cpu.rf_ram.memory[80][5] ),
    .A2(_02614_),
    .ZN(_02620_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06225_ (.A1(_02507_),
    .A2(_02614_),
    .B(_02620_),
    .ZN(_00087_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06226_ (.A1(\u_cpu.rf_ram.memory[80][6] ),
    .A2(_02614_),
    .ZN(_02621_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06227_ (.A1(_02512_),
    .A2(_02614_),
    .B(_02621_),
    .ZN(_00088_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06228_ (.A1(\u_cpu.rf_ram.memory[80][7] ),
    .A2(_02614_),
    .ZN(_02622_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06229_ (.A1(_02517_),
    .A2(_02614_),
    .B(_02622_),
    .ZN(_00089_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _06230_ (.A1(_01386_),
    .A2(_02462_),
    .Z(_02623_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06231_ (.A1(_02522_),
    .A2(_02623_),
    .ZN(_02624_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06232_ (.A1(_02468_),
    .A2(_02624_),
    .ZN(_02625_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06233_ (.A1(_02473_),
    .A2(_02575_),
    .ZN(_02626_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06234_ (.A1(_02625_),
    .A2(_02626_),
    .ZN(_02627_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06235_ (.I(_02627_),
    .Z(_02628_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06236_ (.A1(\u_cpu.rf_ram.memory[78][0] ),
    .A2(_02628_),
    .ZN(_02629_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06237_ (.A1(_02482_),
    .A2(_02628_),
    .B(_02629_),
    .ZN(_00090_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06238_ (.A1(\u_cpu.rf_ram.memory[78][1] ),
    .A2(_02628_),
    .ZN(_02630_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06239_ (.A1(_02487_),
    .A2(_02628_),
    .B(_02630_),
    .ZN(_00091_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06240_ (.A1(\u_cpu.rf_ram.memory[78][2] ),
    .A2(_02628_),
    .ZN(_02631_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06241_ (.A1(_02492_),
    .A2(_02628_),
    .B(_02631_),
    .ZN(_00092_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06242_ (.A1(\u_cpu.rf_ram.memory[78][3] ),
    .A2(_02628_),
    .ZN(_02632_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06243_ (.A1(_02497_),
    .A2(_02628_),
    .B(_02632_),
    .ZN(_00093_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06244_ (.A1(\u_cpu.rf_ram.memory[78][4] ),
    .A2(_02628_),
    .ZN(_02633_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06245_ (.A1(_02502_),
    .A2(_02628_),
    .B(_02633_),
    .ZN(_00094_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06246_ (.A1(\u_cpu.rf_ram.memory[78][5] ),
    .A2(_02628_),
    .ZN(_02634_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06247_ (.A1(_02507_),
    .A2(_02628_),
    .B(_02634_),
    .ZN(_00095_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06248_ (.A1(\u_cpu.rf_ram.memory[78][6] ),
    .A2(_02628_),
    .ZN(_02635_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06249_ (.A1(_02512_),
    .A2(_02628_),
    .B(_02635_),
    .ZN(_00096_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06250_ (.A1(\u_cpu.rf_ram.memory[78][7] ),
    .A2(_02628_),
    .ZN(_02636_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06251_ (.A1(_02517_),
    .A2(_02628_),
    .B(_02636_),
    .ZN(_00097_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06252_ (.A1(_02459_),
    .A2(_02623_),
    .ZN(_02637_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06253_ (.A1(_02468_),
    .A2(_02637_),
    .ZN(_02638_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _06254_ (.A1(\u_cpu.cpu.immdec.imm11_7[2] ),
    .A2(_02526_),
    .A3(_02574_),
    .ZN(_02639_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06255_ (.A1(_02638_),
    .A2(_02639_),
    .ZN(_02640_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06256_ (.I(_02640_),
    .Z(_02641_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06257_ (.A1(\u_cpu.rf_ram.memory[42][0] ),
    .A2(_02641_),
    .ZN(_02642_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06258_ (.A1(_02482_),
    .A2(_02641_),
    .B(_02642_),
    .ZN(_00098_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06259_ (.A1(\u_cpu.rf_ram.memory[42][1] ),
    .A2(_02641_),
    .ZN(_02643_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06260_ (.A1(_02487_),
    .A2(_02641_),
    .B(_02643_),
    .ZN(_00099_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06261_ (.A1(\u_cpu.rf_ram.memory[42][2] ),
    .A2(_02641_),
    .ZN(_02644_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06262_ (.A1(_02492_),
    .A2(_02641_),
    .B(_02644_),
    .ZN(_00100_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06263_ (.A1(\u_cpu.rf_ram.memory[42][3] ),
    .A2(_02641_),
    .ZN(_02645_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06264_ (.A1(_02497_),
    .A2(_02641_),
    .B(_02645_),
    .ZN(_00101_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06265_ (.A1(\u_cpu.rf_ram.memory[42][4] ),
    .A2(_02641_),
    .ZN(_02646_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06266_ (.A1(_02502_),
    .A2(_02641_),
    .B(_02646_),
    .ZN(_00102_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06267_ (.A1(\u_cpu.rf_ram.memory[42][5] ),
    .A2(_02641_),
    .ZN(_02647_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06268_ (.A1(_02507_),
    .A2(_02641_),
    .B(_02647_),
    .ZN(_00103_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06269_ (.A1(\u_cpu.rf_ram.memory[42][6] ),
    .A2(_02641_),
    .ZN(_02648_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06270_ (.A1(_02512_),
    .A2(_02641_),
    .B(_02648_),
    .ZN(_00104_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06271_ (.A1(\u_cpu.rf_ram.memory[42][7] ),
    .A2(_02641_),
    .ZN(_02649_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06272_ (.A1(_02517_),
    .A2(_02641_),
    .B(_02649_),
    .ZN(_00105_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06273_ (.A1(_02625_),
    .A2(_02639_),
    .ZN(_02650_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06274_ (.I(_02650_),
    .Z(_02651_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06275_ (.A1(\u_cpu.rf_ram.memory[46][0] ),
    .A2(_02651_),
    .ZN(_02652_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06276_ (.A1(_02482_),
    .A2(_02651_),
    .B(_02652_),
    .ZN(_00106_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06277_ (.A1(\u_cpu.rf_ram.memory[46][1] ),
    .A2(_02651_),
    .ZN(_02653_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06278_ (.A1(_02487_),
    .A2(_02651_),
    .B(_02653_),
    .ZN(_00107_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06279_ (.A1(\u_cpu.rf_ram.memory[46][2] ),
    .A2(_02651_),
    .ZN(_02654_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06280_ (.A1(_02492_),
    .A2(_02651_),
    .B(_02654_),
    .ZN(_00108_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06281_ (.A1(\u_cpu.rf_ram.memory[46][3] ),
    .A2(_02651_),
    .ZN(_02655_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06282_ (.A1(_02497_),
    .A2(_02651_),
    .B(_02655_),
    .ZN(_00109_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06283_ (.A1(\u_cpu.rf_ram.memory[46][4] ),
    .A2(_02651_),
    .ZN(_02656_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06284_ (.A1(_02502_),
    .A2(_02651_),
    .B(_02656_),
    .ZN(_00110_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06285_ (.A1(\u_cpu.rf_ram.memory[46][5] ),
    .A2(_02651_),
    .ZN(_02657_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06286_ (.A1(_02507_),
    .A2(_02651_),
    .B(_02657_),
    .ZN(_00111_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06287_ (.A1(\u_cpu.rf_ram.memory[46][6] ),
    .A2(_02651_),
    .ZN(_02658_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06288_ (.A1(_02512_),
    .A2(_02651_),
    .B(_02658_),
    .ZN(_00112_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06289_ (.A1(\u_cpu.rf_ram.memory[46][7] ),
    .A2(_02651_),
    .ZN(_02659_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06290_ (.A1(_02517_),
    .A2(_02651_),
    .B(_02659_),
    .ZN(_00113_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06291_ (.A1(_02521_),
    .A2(_02624_),
    .ZN(_02660_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06292_ (.A1(_02639_),
    .A2(_02660_),
    .ZN(_02661_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06293_ (.I(_02661_),
    .Z(_02662_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06294_ (.A1(\u_cpu.rf_ram.memory[45][0] ),
    .A2(_02662_),
    .ZN(_02663_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06295_ (.A1(_02482_),
    .A2(_02662_),
    .B(_02663_),
    .ZN(_00114_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06296_ (.A1(\u_cpu.rf_ram.memory[45][1] ),
    .A2(_02662_),
    .ZN(_02664_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06297_ (.A1(_02487_),
    .A2(_02662_),
    .B(_02664_),
    .ZN(_00115_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06298_ (.A1(\u_cpu.rf_ram.memory[45][2] ),
    .A2(_02662_),
    .ZN(_02665_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06299_ (.A1(_02492_),
    .A2(_02662_),
    .B(_02665_),
    .ZN(_00116_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06300_ (.A1(\u_cpu.rf_ram.memory[45][3] ),
    .A2(_02662_),
    .ZN(_02666_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06301_ (.A1(_02497_),
    .A2(_02662_),
    .B(_02666_),
    .ZN(_00117_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06302_ (.A1(\u_cpu.rf_ram.memory[45][4] ),
    .A2(_02662_),
    .ZN(_02667_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06303_ (.A1(_02502_),
    .A2(_02662_),
    .B(_02667_),
    .ZN(_00118_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06304_ (.A1(\u_cpu.rf_ram.memory[45][5] ),
    .A2(_02662_),
    .ZN(_02668_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06305_ (.A1(_02507_),
    .A2(_02662_),
    .B(_02668_),
    .ZN(_00119_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06306_ (.A1(\u_cpu.rf_ram.memory[45][6] ),
    .A2(_02662_),
    .ZN(_02669_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06307_ (.A1(_02512_),
    .A2(_02662_),
    .B(_02669_),
    .ZN(_00120_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06308_ (.A1(\u_cpu.rf_ram.memory[45][7] ),
    .A2(_02662_),
    .ZN(_02670_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06309_ (.A1(_02517_),
    .A2(_02662_),
    .B(_02670_),
    .ZN(_00121_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06310_ (.A1(_02560_),
    .A2(_02624_),
    .ZN(_02671_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06311_ (.A1(_02639_),
    .A2(_02671_),
    .ZN(_02672_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06312_ (.I(_02672_),
    .Z(_02673_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06313_ (.A1(\u_cpu.rf_ram.memory[44][0] ),
    .A2(_02673_),
    .ZN(_02674_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06314_ (.A1(_02482_),
    .A2(_02673_),
    .B(_02674_),
    .ZN(_00122_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06315_ (.A1(\u_cpu.rf_ram.memory[44][1] ),
    .A2(_02673_),
    .ZN(_02675_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06316_ (.A1(_02487_),
    .A2(_02673_),
    .B(_02675_),
    .ZN(_00123_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06317_ (.A1(\u_cpu.rf_ram.memory[44][2] ),
    .A2(_02673_),
    .ZN(_02676_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06318_ (.A1(_02492_),
    .A2(_02673_),
    .B(_02676_),
    .ZN(_00124_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06319_ (.A1(\u_cpu.rf_ram.memory[44][3] ),
    .A2(_02673_),
    .ZN(_02677_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06320_ (.A1(_02497_),
    .A2(_02673_),
    .B(_02677_),
    .ZN(_00125_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06321_ (.A1(\u_cpu.rf_ram.memory[44][4] ),
    .A2(_02673_),
    .ZN(_02678_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06322_ (.A1(_02502_),
    .A2(_02673_),
    .B(_02678_),
    .ZN(_00126_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06323_ (.A1(\u_cpu.rf_ram.memory[44][5] ),
    .A2(_02673_),
    .ZN(_02679_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06324_ (.A1(_02507_),
    .A2(_02673_),
    .B(_02679_),
    .ZN(_00127_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06325_ (.A1(\u_cpu.rf_ram.memory[44][6] ),
    .A2(_02673_),
    .ZN(_02680_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06326_ (.A1(_02512_),
    .A2(_02673_),
    .B(_02680_),
    .ZN(_00128_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06327_ (.A1(\u_cpu.rf_ram.memory[44][7] ),
    .A2(_02673_),
    .ZN(_02681_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06328_ (.A1(_02517_),
    .A2(_02673_),
    .B(_02681_),
    .ZN(_00129_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06329_ (.A1(_02464_),
    .A2(_02601_),
    .ZN(_02682_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06330_ (.A1(\u_cpu.cpu.immdec.imm11_7[2] ),
    .A2(\u_cpu.cpu.immdec.imm11_7[3] ),
    .A3(_02457_),
    .ZN(_02683_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06331_ (.A1(_02526_),
    .A2(_02683_),
    .ZN(_02684_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06332_ (.A1(_02682_),
    .A2(_02684_),
    .ZN(_02685_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06333_ (.I(_02685_),
    .Z(_02686_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06334_ (.A1(\u_cpu.rf_ram.memory[51][0] ),
    .A2(_02686_),
    .ZN(_02687_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06335_ (.A1(_02482_),
    .A2(_02686_),
    .B(_02687_),
    .ZN(_00130_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06336_ (.A1(\u_cpu.rf_ram.memory[51][1] ),
    .A2(_02686_),
    .ZN(_02688_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06337_ (.A1(_02487_),
    .A2(_02686_),
    .B(_02688_),
    .ZN(_00131_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06338_ (.A1(\u_cpu.rf_ram.memory[51][2] ),
    .A2(_02686_),
    .ZN(_02689_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06339_ (.A1(_02492_),
    .A2(_02686_),
    .B(_02689_),
    .ZN(_00132_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06340_ (.A1(\u_cpu.rf_ram.memory[51][3] ),
    .A2(_02686_),
    .ZN(_02690_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06341_ (.A1(_02497_),
    .A2(_02686_),
    .B(_02690_),
    .ZN(_00133_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06342_ (.A1(\u_cpu.rf_ram.memory[51][4] ),
    .A2(_02686_),
    .ZN(_02691_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06343_ (.A1(_02502_),
    .A2(_02686_),
    .B(_02691_),
    .ZN(_00134_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06344_ (.A1(\u_cpu.rf_ram.memory[51][5] ),
    .A2(_02686_),
    .ZN(_02692_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06345_ (.A1(_02507_),
    .A2(_02686_),
    .B(_02692_),
    .ZN(_00135_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06346_ (.A1(\u_cpu.rf_ram.memory[51][6] ),
    .A2(_02686_),
    .ZN(_02693_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06347_ (.A1(_02512_),
    .A2(_02686_),
    .B(_02693_),
    .ZN(_00136_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06348_ (.A1(\u_cpu.rf_ram.memory[51][7] ),
    .A2(_02686_),
    .ZN(_02694_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06349_ (.A1(_02517_),
    .A2(_02686_),
    .B(_02694_),
    .ZN(_00137_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06350_ (.A1(_02521_),
    .A2(_02637_),
    .ZN(_02695_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06351_ (.A1(_02639_),
    .A2(_02695_),
    .ZN(_02696_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06352_ (.I(_02696_),
    .Z(_02697_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06353_ (.A1(\u_cpu.rf_ram.memory[41][0] ),
    .A2(_02697_),
    .ZN(_02698_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06354_ (.A1(_02482_),
    .A2(_02697_),
    .B(_02698_),
    .ZN(_00138_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06355_ (.A1(\u_cpu.rf_ram.memory[41][1] ),
    .A2(_02697_),
    .ZN(_02699_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06356_ (.A1(_02487_),
    .A2(_02697_),
    .B(_02699_),
    .ZN(_00139_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06357_ (.A1(\u_cpu.rf_ram.memory[41][2] ),
    .A2(_02697_),
    .ZN(_02700_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06358_ (.A1(_02492_),
    .A2(_02697_),
    .B(_02700_),
    .ZN(_00140_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06359_ (.A1(\u_cpu.rf_ram.memory[41][3] ),
    .A2(_02697_),
    .ZN(_02701_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06360_ (.A1(_02497_),
    .A2(_02697_),
    .B(_02701_),
    .ZN(_00141_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06361_ (.A1(\u_cpu.rf_ram.memory[41][4] ),
    .A2(_02697_),
    .ZN(_02702_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06362_ (.A1(_02502_),
    .A2(_02697_),
    .B(_02702_),
    .ZN(_00142_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06363_ (.A1(\u_cpu.rf_ram.memory[41][5] ),
    .A2(_02697_),
    .ZN(_02703_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06364_ (.A1(_02507_),
    .A2(_02697_),
    .B(_02703_),
    .ZN(_00143_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06365_ (.A1(\u_cpu.rf_ram.memory[41][6] ),
    .A2(_02697_),
    .ZN(_02704_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06366_ (.A1(_02512_),
    .A2(_02697_),
    .B(_02704_),
    .ZN(_00144_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06367_ (.A1(\u_cpu.rf_ram.memory[41][7] ),
    .A2(_02697_),
    .ZN(_02705_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06368_ (.A1(_02517_),
    .A2(_02697_),
    .B(_02705_),
    .ZN(_00145_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06369_ (.A1(_02601_),
    .A2(_02637_),
    .ZN(_02706_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06370_ (.A1(_02639_),
    .A2(_02706_),
    .ZN(_02707_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06371_ (.I(_02707_),
    .Z(_02708_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06372_ (.A1(\u_cpu.rf_ram.memory[43][0] ),
    .A2(_02708_),
    .ZN(_02709_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06373_ (.A1(_02482_),
    .A2(_02708_),
    .B(_02709_),
    .ZN(_00146_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06374_ (.A1(\u_cpu.rf_ram.memory[43][1] ),
    .A2(_02708_),
    .ZN(_02710_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06375_ (.A1(_02487_),
    .A2(_02708_),
    .B(_02710_),
    .ZN(_00147_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06376_ (.A1(\u_cpu.rf_ram.memory[43][2] ),
    .A2(_02708_),
    .ZN(_02711_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06377_ (.A1(_02492_),
    .A2(_02708_),
    .B(_02711_),
    .ZN(_00148_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06378_ (.A1(\u_cpu.rf_ram.memory[43][3] ),
    .A2(_02708_),
    .ZN(_02712_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06379_ (.A1(_02497_),
    .A2(_02708_),
    .B(_02712_),
    .ZN(_00149_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06380_ (.A1(\u_cpu.rf_ram.memory[43][4] ),
    .A2(_02708_),
    .ZN(_02713_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06381_ (.A1(_02502_),
    .A2(_02708_),
    .B(_02713_),
    .ZN(_00150_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06382_ (.A1(\u_cpu.rf_ram.memory[43][5] ),
    .A2(_02708_),
    .ZN(_02714_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06383_ (.A1(_02507_),
    .A2(_02708_),
    .B(_02714_),
    .ZN(_00151_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06384_ (.A1(\u_cpu.rf_ram.memory[43][6] ),
    .A2(_02708_),
    .ZN(_02715_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06385_ (.A1(_02512_),
    .A2(_02708_),
    .B(_02715_),
    .ZN(_00152_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06386_ (.A1(\u_cpu.rf_ram.memory[43][7] ),
    .A2(_02708_),
    .ZN(_02716_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06387_ (.A1(_02517_),
    .A2(_02708_),
    .B(_02716_),
    .ZN(_00153_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06388_ (.A1(_02612_),
    .A2(_02684_),
    .ZN(_02717_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06389_ (.I(_02717_),
    .Z(_02718_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06390_ (.A1(\u_cpu.rf_ram.memory[48][0] ),
    .A2(_02718_),
    .ZN(_02719_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06391_ (.A1(_02482_),
    .A2(_02718_),
    .B(_02719_),
    .ZN(_00154_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06392_ (.A1(\u_cpu.rf_ram.memory[48][1] ),
    .A2(_02718_),
    .ZN(_02720_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06393_ (.A1(_02487_),
    .A2(_02718_),
    .B(_02720_),
    .ZN(_00155_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06394_ (.A1(\u_cpu.rf_ram.memory[48][2] ),
    .A2(_02718_),
    .ZN(_02721_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06395_ (.A1(_02492_),
    .A2(_02718_),
    .B(_02721_),
    .ZN(_00156_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06396_ (.A1(\u_cpu.rf_ram.memory[48][3] ),
    .A2(_02718_),
    .ZN(_02722_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06397_ (.A1(_02497_),
    .A2(_02718_),
    .B(_02722_),
    .ZN(_00157_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06398_ (.A1(\u_cpu.rf_ram.memory[48][4] ),
    .A2(_02718_),
    .ZN(_02723_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06399_ (.A1(_02502_),
    .A2(_02718_),
    .B(_02723_),
    .ZN(_00158_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06400_ (.A1(\u_cpu.rf_ram.memory[48][5] ),
    .A2(_02718_),
    .ZN(_02724_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06401_ (.A1(_02507_),
    .A2(_02718_),
    .B(_02724_),
    .ZN(_00159_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06402_ (.A1(\u_cpu.rf_ram.memory[48][6] ),
    .A2(_02718_),
    .ZN(_02725_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06403_ (.A1(_02512_),
    .A2(_02718_),
    .B(_02725_),
    .ZN(_00160_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06404_ (.A1(\u_cpu.rf_ram.memory[48][7] ),
    .A2(_02718_),
    .ZN(_02726_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06405_ (.A1(_02517_),
    .A2(_02718_),
    .B(_02726_),
    .ZN(_00161_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06406_ (.A1(_02601_),
    .A2(_02624_),
    .ZN(_02727_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06407_ (.A1(_02639_),
    .A2(_02727_),
    .ZN(_02728_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06408_ (.I(_02728_),
    .Z(_02729_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06409_ (.A1(\u_cpu.rf_ram.memory[47][0] ),
    .A2(_02729_),
    .ZN(_02730_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06410_ (.A1(_02482_),
    .A2(_02729_),
    .B(_02730_),
    .ZN(_00162_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06411_ (.A1(\u_cpu.rf_ram.memory[47][1] ),
    .A2(_02729_),
    .ZN(_02731_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06412_ (.A1(_02487_),
    .A2(_02729_),
    .B(_02731_),
    .ZN(_00163_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06413_ (.A1(\u_cpu.rf_ram.memory[47][2] ),
    .A2(_02729_),
    .ZN(_02732_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06414_ (.A1(_02492_),
    .A2(_02729_),
    .B(_02732_),
    .ZN(_00164_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06415_ (.A1(\u_cpu.rf_ram.memory[47][3] ),
    .A2(_02729_),
    .ZN(_02733_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06416_ (.A1(_02497_),
    .A2(_02729_),
    .B(_02733_),
    .ZN(_00165_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06417_ (.A1(\u_cpu.rf_ram.memory[47][4] ),
    .A2(_02729_),
    .ZN(_02734_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06418_ (.A1(_02502_),
    .A2(_02729_),
    .B(_02734_),
    .ZN(_00166_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06419_ (.A1(\u_cpu.rf_ram.memory[47][5] ),
    .A2(_02729_),
    .ZN(_02735_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06420_ (.A1(_02507_),
    .A2(_02729_),
    .B(_02735_),
    .ZN(_00167_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06421_ (.A1(\u_cpu.rf_ram.memory[47][6] ),
    .A2(_02729_),
    .ZN(_02736_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06422_ (.A1(_02512_),
    .A2(_02729_),
    .B(_02736_),
    .ZN(_00168_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06423_ (.A1(\u_cpu.rf_ram.memory[47][7] ),
    .A2(_02729_),
    .ZN(_02737_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06424_ (.A1(_02517_),
    .A2(_02729_),
    .B(_02737_),
    .ZN(_00169_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06425_ (.I(_02481_),
    .Z(_02738_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06426_ (.A1(_02469_),
    .A2(_02684_),
    .ZN(_02739_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06427_ (.I(_02739_),
    .Z(_02740_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06428_ (.A1(\u_cpu.rf_ram.memory[50][0] ),
    .A2(_02740_),
    .ZN(_02741_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06429_ (.A1(_02738_),
    .A2(_02740_),
    .B(_02741_),
    .ZN(_00170_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06430_ (.I(_02486_),
    .Z(_02742_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06431_ (.A1(\u_cpu.rf_ram.memory[50][1] ),
    .A2(_02740_),
    .ZN(_02743_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06432_ (.A1(_02742_),
    .A2(_02740_),
    .B(_02743_),
    .ZN(_00171_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06433_ (.I(_02491_),
    .Z(_02744_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06434_ (.A1(\u_cpu.rf_ram.memory[50][2] ),
    .A2(_02740_),
    .ZN(_02745_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06435_ (.A1(_02744_),
    .A2(_02740_),
    .B(_02745_),
    .ZN(_00172_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06436_ (.I(_02496_),
    .Z(_02746_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06437_ (.A1(\u_cpu.rf_ram.memory[50][3] ),
    .A2(_02740_),
    .ZN(_02747_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06438_ (.A1(_02746_),
    .A2(_02740_),
    .B(_02747_),
    .ZN(_00173_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06439_ (.I(_02501_),
    .Z(_02748_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06440_ (.A1(\u_cpu.rf_ram.memory[50][4] ),
    .A2(_02740_),
    .ZN(_02749_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06441_ (.A1(_02748_),
    .A2(_02740_),
    .B(_02749_),
    .ZN(_00174_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06442_ (.I(_02506_),
    .Z(_02750_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06443_ (.A1(\u_cpu.rf_ram.memory[50][5] ),
    .A2(_02740_),
    .ZN(_02751_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06444_ (.A1(_02750_),
    .A2(_02740_),
    .B(_02751_),
    .ZN(_00175_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06445_ (.I(_02511_),
    .Z(_02752_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06446_ (.A1(\u_cpu.rf_ram.memory[50][6] ),
    .A2(_02740_),
    .ZN(_02753_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06447_ (.A1(_02752_),
    .A2(_02740_),
    .B(_02753_),
    .ZN(_00176_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06448_ (.I(_02516_),
    .Z(_02754_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06449_ (.A1(\u_cpu.rf_ram.memory[50][7] ),
    .A2(_02740_),
    .ZN(_02755_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06450_ (.A1(_02754_),
    .A2(_02740_),
    .B(_02755_),
    .ZN(_00177_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06451_ (.A1(_02561_),
    .A2(_02577_),
    .ZN(_02756_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06452_ (.I0(_02573_),
    .I1(\u_cpu.rf_ram.memory[4][0] ),
    .S(_02756_),
    .Z(_02757_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06453_ (.I(_02757_),
    .Z(_00178_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06454_ (.I0(_02581_),
    .I1(\u_cpu.rf_ram.memory[4][1] ),
    .S(_02756_),
    .Z(_02758_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06455_ (.I(_02758_),
    .Z(_00179_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06456_ (.I0(_02584_),
    .I1(\u_cpu.rf_ram.memory[4][2] ),
    .S(_02756_),
    .Z(_02759_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06457_ (.I(_02759_),
    .Z(_00180_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06458_ (.I0(_02587_),
    .I1(\u_cpu.rf_ram.memory[4][3] ),
    .S(_02756_),
    .Z(_02760_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06459_ (.I(_02760_),
    .Z(_00181_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06460_ (.I0(_02590_),
    .I1(\u_cpu.rf_ram.memory[4][4] ),
    .S(_02756_),
    .Z(_02761_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06461_ (.I(_02761_),
    .Z(_00182_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06462_ (.I0(_02593_),
    .I1(\u_cpu.rf_ram.memory[4][5] ),
    .S(_02756_),
    .Z(_02762_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06463_ (.I(_02762_),
    .Z(_00183_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06464_ (.I0(_02596_),
    .I1(\u_cpu.rf_ram.memory[4][6] ),
    .S(_02756_),
    .Z(_02763_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06465_ (.I(_02763_),
    .Z(_00184_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06466_ (.I0(_02599_),
    .I1(\u_cpu.rf_ram.memory[4][7] ),
    .S(_02756_),
    .Z(_02764_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06467_ (.I(_02764_),
    .Z(_00185_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _06468_ (.I(_01435_),
    .ZN(_02765_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06469_ (.A1(\u_arbiter.i_wb_cpu_ack ),
    .A2(_01431_),
    .ZN(_02766_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06470_ (.A1(_02765_),
    .A2(\u_arbiter.i_wb_cpu_ibus_adr[1] ),
    .B(_02766_),
    .ZN(_02767_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06471_ (.I(_02767_),
    .Z(_02768_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06472_ (.A1(\u_cpu.cpu.state.genblk1.misalign_trap_sync_r ),
    .A2(\u_cpu.cpu.state.stage_two_req ),
    .B(_02768_),
    .ZN(_02769_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06473_ (.A1(_01428_),
    .A2(_02769_),
    .ZN(_00186_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06474_ (.A1(_02311_),
    .A2(_02448_),
    .B(_02367_),
    .ZN(_02770_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06475_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[6] ),
    .A2(_02770_),
    .ZN(_02771_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06476_ (.A1(_01372_),
    .A2(_02332_),
    .ZN(_02772_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06477_ (.A1(_02447_),
    .A2(_02365_),
    .Z(_02773_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06478_ (.A1(_02772_),
    .A2(_02773_),
    .ZN(_02774_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _06479_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[0] ),
    .A2(\u_arbiter.i_wb_cpu_dbus_dat[1] ),
    .A3(\u_arbiter.i_wb_cpu_dbus_dat[2] ),
    .A4(\u_arbiter.i_wb_cpu_dbus_dat[3] ),
    .Z(_02775_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06480_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[4] ),
    .A2(_02775_),
    .ZN(_02776_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06481_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[5] ),
    .A2(_02776_),
    .Z(_02777_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06482_ (.A1(_02774_),
    .A2(_02777_),
    .ZN(_02778_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06483_ (.A1(_02771_),
    .A2(_02778_),
    .ZN(_02779_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _06484_ (.A1(_01408_),
    .A2(_01370_),
    .A3(_02779_),
    .ZN(_02780_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06485_ (.A1(\u_arbiter.i_wb_cpu_ack ),
    .A2(_01442_),
    .ZN(_02781_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _06486_ (.A1(_01373_),
    .A2(_02780_),
    .B(_02781_),
    .C(_01375_),
    .ZN(_02782_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _06487_ (.A1(\u_cpu.cpu.state.init_done ),
    .A2(_01385_),
    .A3(_02433_),
    .A4(_02782_),
    .ZN(_02783_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06488_ (.A1(_02769_),
    .A2(_02783_),
    .ZN(_02784_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06489_ (.A1(\u_cpu.rf_ram_if.rcnt[0] ),
    .A2(_02784_),
    .ZN(_00187_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _06490_ (.A1(\u_cpu.rf_ram_if.rcnt[2] ),
    .A2(\u_cpu.rf_ram_if.rcnt[1] ),
    .A3(\u_cpu.rf_ram_if.rcnt[0] ),
    .Z(_02785_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _06491_ (.A1(_02465_),
    .A2(_02784_),
    .A3(_02785_),
    .ZN(_00188_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06492_ (.A1(_01680_),
    .A2(_02785_),
    .ZN(_02786_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _06493_ (.A1(_01680_),
    .A2(_02785_),
    .Z(_02787_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _06494_ (.A1(_02769_),
    .A2(_02783_),
    .A3(_02786_),
    .A4(_02787_),
    .Z(_02788_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06495_ (.I(_02788_),
    .Z(_00189_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06496_ (.A1(_01681_),
    .A2(_02786_),
    .Z(_02789_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06497_ (.A1(_02784_),
    .A2(_02789_),
    .ZN(_00190_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06498_ (.A1(_02528_),
    .A2(_02612_),
    .ZN(_02790_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06499_ (.I(_02790_),
    .Z(_02791_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06500_ (.A1(\u_cpu.rf_ram.memory[16][0] ),
    .A2(_02791_),
    .ZN(_02792_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06501_ (.A1(_02738_),
    .A2(_02791_),
    .B(_02792_),
    .ZN(_00191_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06502_ (.A1(\u_cpu.rf_ram.memory[16][1] ),
    .A2(_02791_),
    .ZN(_02793_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06503_ (.A1(_02742_),
    .A2(_02791_),
    .B(_02793_),
    .ZN(_00192_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06504_ (.A1(\u_cpu.rf_ram.memory[16][2] ),
    .A2(_02791_),
    .ZN(_02794_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06505_ (.A1(_02744_),
    .A2(_02791_),
    .B(_02794_),
    .ZN(_00193_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06506_ (.A1(\u_cpu.rf_ram.memory[16][3] ),
    .A2(_02791_),
    .ZN(_02795_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06507_ (.A1(_02746_),
    .A2(_02791_),
    .B(_02795_),
    .ZN(_00194_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06508_ (.A1(\u_cpu.rf_ram.memory[16][4] ),
    .A2(_02791_),
    .ZN(_02796_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06509_ (.A1(_02748_),
    .A2(_02791_),
    .B(_02796_),
    .ZN(_00195_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06510_ (.A1(\u_cpu.rf_ram.memory[16][5] ),
    .A2(_02791_),
    .ZN(_02797_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06511_ (.A1(_02750_),
    .A2(_02791_),
    .B(_02797_),
    .ZN(_00196_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06512_ (.A1(\u_cpu.rf_ram.memory[16][6] ),
    .A2(_02791_),
    .ZN(_02798_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06513_ (.A1(_02752_),
    .A2(_02791_),
    .B(_02798_),
    .ZN(_00197_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06514_ (.A1(\u_cpu.rf_ram.memory[16][7] ),
    .A2(_02791_),
    .ZN(_02799_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06515_ (.A1(_02754_),
    .A2(_02791_),
    .B(_02799_),
    .ZN(_00198_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06516_ (.A1(_02528_),
    .A2(_02539_),
    .ZN(_02800_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06517_ (.I(_02800_),
    .Z(_02801_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06518_ (.A1(\u_cpu.rf_ram.memory[17][0] ),
    .A2(_02801_),
    .ZN(_02802_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06519_ (.A1(_02738_),
    .A2(_02801_),
    .B(_02802_),
    .ZN(_00199_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06520_ (.A1(\u_cpu.rf_ram.memory[17][1] ),
    .A2(_02801_),
    .ZN(_02803_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06521_ (.A1(_02742_),
    .A2(_02801_),
    .B(_02803_),
    .ZN(_00200_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06522_ (.A1(\u_cpu.rf_ram.memory[17][2] ),
    .A2(_02801_),
    .ZN(_02804_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06523_ (.A1(_02744_),
    .A2(_02801_),
    .B(_02804_),
    .ZN(_00201_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06524_ (.A1(\u_cpu.rf_ram.memory[17][3] ),
    .A2(_02801_),
    .ZN(_02805_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06525_ (.A1(_02746_),
    .A2(_02801_),
    .B(_02805_),
    .ZN(_00202_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06526_ (.A1(\u_cpu.rf_ram.memory[17][4] ),
    .A2(_02801_),
    .ZN(_02806_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06527_ (.A1(_02748_),
    .A2(_02801_),
    .B(_02806_),
    .ZN(_00203_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06528_ (.A1(\u_cpu.rf_ram.memory[17][5] ),
    .A2(_02801_),
    .ZN(_02807_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06529_ (.A1(_02750_),
    .A2(_02801_),
    .B(_02807_),
    .ZN(_00204_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06530_ (.A1(\u_cpu.rf_ram.memory[17][6] ),
    .A2(_02801_),
    .ZN(_02808_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06531_ (.A1(_02752_),
    .A2(_02801_),
    .B(_02808_),
    .ZN(_00205_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06532_ (.A1(\u_cpu.rf_ram.memory[17][7] ),
    .A2(_02801_),
    .ZN(_02809_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06533_ (.A1(_02754_),
    .A2(_02801_),
    .B(_02809_),
    .ZN(_00206_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06534_ (.A1(_02560_),
    .A2(_02637_),
    .ZN(_02810_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06535_ (.A1(_02639_),
    .A2(_02810_),
    .ZN(_02811_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06536_ (.I(_02811_),
    .Z(_02812_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06537_ (.A1(\u_cpu.rf_ram.memory[40][0] ),
    .A2(_02812_),
    .ZN(_02813_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06538_ (.A1(_02738_),
    .A2(_02812_),
    .B(_02813_),
    .ZN(_00207_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06539_ (.A1(\u_cpu.rf_ram.memory[40][1] ),
    .A2(_02812_),
    .ZN(_02814_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06540_ (.A1(_02742_),
    .A2(_02812_),
    .B(_02814_),
    .ZN(_00208_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06541_ (.A1(\u_cpu.rf_ram.memory[40][2] ),
    .A2(_02812_),
    .ZN(_02815_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06542_ (.A1(_02744_),
    .A2(_02812_),
    .B(_02815_),
    .ZN(_00209_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06543_ (.A1(\u_cpu.rf_ram.memory[40][3] ),
    .A2(_02812_),
    .ZN(_02816_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06544_ (.A1(_02746_),
    .A2(_02812_),
    .B(_02816_),
    .ZN(_00210_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06545_ (.A1(\u_cpu.rf_ram.memory[40][4] ),
    .A2(_02812_),
    .ZN(_02817_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06546_ (.A1(_02748_),
    .A2(_02812_),
    .B(_02817_),
    .ZN(_00211_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06547_ (.A1(\u_cpu.rf_ram.memory[40][5] ),
    .A2(_02812_),
    .ZN(_02818_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06548_ (.A1(_02750_),
    .A2(_02812_),
    .B(_02818_),
    .ZN(_00212_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06549_ (.A1(\u_cpu.rf_ram.memory[40][6] ),
    .A2(_02812_),
    .ZN(_02819_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06550_ (.A1(_02752_),
    .A2(_02812_),
    .B(_02819_),
    .ZN(_00213_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06551_ (.A1(\u_cpu.rf_ram.memory[40][7] ),
    .A2(_02812_),
    .ZN(_02820_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06552_ (.A1(_02754_),
    .A2(_02812_),
    .B(_02820_),
    .ZN(_00214_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06553_ (.A1(_02473_),
    .A2(_02683_),
    .ZN(_02821_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06554_ (.A1(_02602_),
    .A2(_02821_),
    .ZN(_02822_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06555_ (.I(_02822_),
    .Z(_02823_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06556_ (.A1(\u_cpu.rf_ram.memory[119][0] ),
    .A2(_02823_),
    .ZN(_02824_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06557_ (.A1(_02738_),
    .A2(_02823_),
    .B(_02824_),
    .ZN(_00215_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06558_ (.A1(\u_cpu.rf_ram.memory[119][1] ),
    .A2(_02823_),
    .ZN(_02825_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06559_ (.A1(_02742_),
    .A2(_02823_),
    .B(_02825_),
    .ZN(_00216_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06560_ (.A1(\u_cpu.rf_ram.memory[119][2] ),
    .A2(_02823_),
    .ZN(_02826_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06561_ (.A1(_02744_),
    .A2(_02823_),
    .B(_02826_),
    .ZN(_00217_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06562_ (.A1(\u_cpu.rf_ram.memory[119][3] ),
    .A2(_02823_),
    .ZN(_02827_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06563_ (.A1(_02746_),
    .A2(_02823_),
    .B(_02827_),
    .ZN(_00218_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06564_ (.A1(\u_cpu.rf_ram.memory[119][4] ),
    .A2(_02823_),
    .ZN(_02828_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06565_ (.A1(_02748_),
    .A2(_02823_),
    .B(_02828_),
    .ZN(_00219_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06566_ (.A1(\u_cpu.rf_ram.memory[119][5] ),
    .A2(_02823_),
    .ZN(_02829_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06567_ (.A1(_02750_),
    .A2(_02823_),
    .B(_02829_),
    .ZN(_00220_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06568_ (.A1(\u_cpu.rf_ram.memory[119][6] ),
    .A2(_02823_),
    .ZN(_02830_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06569_ (.A1(_02752_),
    .A2(_02823_),
    .B(_02830_),
    .ZN(_00221_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06570_ (.A1(\u_cpu.rf_ram.memory[119][7] ),
    .A2(_02823_),
    .ZN(_02831_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06571_ (.A1(_02754_),
    .A2(_02823_),
    .B(_02831_),
    .ZN(_00222_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06572_ (.A1(_02457_),
    .A2(_02471_),
    .ZN(_02832_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06573_ (.A1(_02539_),
    .A2(_02832_),
    .ZN(_02833_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06574_ (.I(_02833_),
    .Z(_02834_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06575_ (.A1(\u_cpu.rf_ram.memory[129][0] ),
    .A2(_02834_),
    .ZN(_02835_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06576_ (.A1(_02738_),
    .A2(_02834_),
    .B(_02835_),
    .ZN(_00223_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06577_ (.A1(\u_cpu.rf_ram.memory[129][1] ),
    .A2(_02834_),
    .ZN(_02836_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06578_ (.A1(_02742_),
    .A2(_02834_),
    .B(_02836_),
    .ZN(_00224_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06579_ (.A1(\u_cpu.rf_ram.memory[129][2] ),
    .A2(_02834_),
    .ZN(_02837_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06580_ (.A1(_02744_),
    .A2(_02834_),
    .B(_02837_),
    .ZN(_00225_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06581_ (.A1(\u_cpu.rf_ram.memory[129][3] ),
    .A2(_02834_),
    .ZN(_02838_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06582_ (.A1(_02746_),
    .A2(_02834_),
    .B(_02838_),
    .ZN(_00226_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06583_ (.A1(\u_cpu.rf_ram.memory[129][4] ),
    .A2(_02834_),
    .ZN(_02839_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06584_ (.A1(_02748_),
    .A2(_02834_),
    .B(_02839_),
    .ZN(_00227_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06585_ (.A1(\u_cpu.rf_ram.memory[129][5] ),
    .A2(_02834_),
    .ZN(_02840_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06586_ (.A1(_02750_),
    .A2(_02834_),
    .B(_02840_),
    .ZN(_00228_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06587_ (.A1(\u_cpu.rf_ram.memory[129][6] ),
    .A2(_02834_),
    .ZN(_02841_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06588_ (.A1(_02752_),
    .A2(_02834_),
    .B(_02841_),
    .ZN(_00229_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06589_ (.A1(\u_cpu.rf_ram.memory[129][7] ),
    .A2(_02834_),
    .ZN(_02842_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06590_ (.A1(_02754_),
    .A2(_02834_),
    .B(_02842_),
    .ZN(_00230_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06591_ (.A1(_02706_),
    .A2(_02832_),
    .ZN(_02843_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06592_ (.I(_02843_),
    .Z(_02844_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06593_ (.A1(\u_cpu.rf_ram.memory[139][0] ),
    .A2(_02844_),
    .ZN(_02845_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06594_ (.A1(_02738_),
    .A2(_02844_),
    .B(_02845_),
    .ZN(_00231_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06595_ (.A1(\u_cpu.rf_ram.memory[139][1] ),
    .A2(_02844_),
    .ZN(_02846_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06596_ (.A1(_02742_),
    .A2(_02844_),
    .B(_02846_),
    .ZN(_00232_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06597_ (.A1(\u_cpu.rf_ram.memory[139][2] ),
    .A2(_02844_),
    .ZN(_02847_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06598_ (.A1(_02744_),
    .A2(_02844_),
    .B(_02847_),
    .ZN(_00233_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06599_ (.A1(\u_cpu.rf_ram.memory[139][3] ),
    .A2(_02844_),
    .ZN(_02848_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06600_ (.A1(_02746_),
    .A2(_02844_),
    .B(_02848_),
    .ZN(_00234_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06601_ (.A1(\u_cpu.rf_ram.memory[139][4] ),
    .A2(_02844_),
    .ZN(_02849_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06602_ (.A1(_02748_),
    .A2(_02844_),
    .B(_02849_),
    .ZN(_00235_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06603_ (.A1(\u_cpu.rf_ram.memory[139][5] ),
    .A2(_02844_),
    .ZN(_02850_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06604_ (.A1(_02750_),
    .A2(_02844_),
    .B(_02850_),
    .ZN(_00236_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06605_ (.A1(\u_cpu.rf_ram.memory[139][6] ),
    .A2(_02844_),
    .ZN(_02851_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06606_ (.A1(_02752_),
    .A2(_02844_),
    .B(_02851_),
    .ZN(_00237_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06607_ (.A1(\u_cpu.rf_ram.memory[139][7] ),
    .A2(_02844_),
    .ZN(_02852_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06608_ (.A1(_02754_),
    .A2(_02844_),
    .B(_02852_),
    .ZN(_00238_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06609_ (.A1(_02626_),
    .A2(_02660_),
    .ZN(_02853_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06610_ (.I(_02853_),
    .Z(_02854_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06611_ (.A1(\u_cpu.rf_ram.memory[77][0] ),
    .A2(_02854_),
    .ZN(_02855_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06612_ (.A1(_02738_),
    .A2(_02854_),
    .B(_02855_),
    .ZN(_00239_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06613_ (.A1(\u_cpu.rf_ram.memory[77][1] ),
    .A2(_02854_),
    .ZN(_02856_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06614_ (.A1(_02742_),
    .A2(_02854_),
    .B(_02856_),
    .ZN(_00240_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06615_ (.A1(\u_cpu.rf_ram.memory[77][2] ),
    .A2(_02854_),
    .ZN(_02857_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06616_ (.A1(_02744_),
    .A2(_02854_),
    .B(_02857_),
    .ZN(_00241_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06617_ (.A1(\u_cpu.rf_ram.memory[77][3] ),
    .A2(_02854_),
    .ZN(_02858_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06618_ (.A1(_02746_),
    .A2(_02854_),
    .B(_02858_),
    .ZN(_00242_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06619_ (.A1(\u_cpu.rf_ram.memory[77][4] ),
    .A2(_02854_),
    .ZN(_02859_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06620_ (.A1(_02748_),
    .A2(_02854_),
    .B(_02859_),
    .ZN(_00243_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06621_ (.A1(\u_cpu.rf_ram.memory[77][5] ),
    .A2(_02854_),
    .ZN(_02860_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06622_ (.A1(_02750_),
    .A2(_02854_),
    .B(_02860_),
    .ZN(_00244_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06623_ (.A1(\u_cpu.rf_ram.memory[77][6] ),
    .A2(_02854_),
    .ZN(_02861_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06624_ (.A1(_02752_),
    .A2(_02854_),
    .B(_02861_),
    .ZN(_00245_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06625_ (.A1(\u_cpu.rf_ram.memory[77][7] ),
    .A2(_02854_),
    .ZN(_02862_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06626_ (.A1(_02754_),
    .A2(_02854_),
    .B(_02862_),
    .ZN(_00246_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06627_ (.A1(_02626_),
    .A2(_02638_),
    .ZN(_02863_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06628_ (.I(_02863_),
    .Z(_02864_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06629_ (.A1(\u_cpu.rf_ram.memory[74][0] ),
    .A2(_02864_),
    .ZN(_02865_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06630_ (.A1(_02738_),
    .A2(_02864_),
    .B(_02865_),
    .ZN(_00247_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06631_ (.A1(\u_cpu.rf_ram.memory[74][1] ),
    .A2(_02864_),
    .ZN(_02866_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06632_ (.A1(_02742_),
    .A2(_02864_),
    .B(_02866_),
    .ZN(_00248_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06633_ (.A1(\u_cpu.rf_ram.memory[74][2] ),
    .A2(_02864_),
    .ZN(_02867_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06634_ (.A1(_02744_),
    .A2(_02864_),
    .B(_02867_),
    .ZN(_00249_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06635_ (.A1(\u_cpu.rf_ram.memory[74][3] ),
    .A2(_02864_),
    .ZN(_02868_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06636_ (.A1(_02746_),
    .A2(_02864_),
    .B(_02868_),
    .ZN(_00250_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06637_ (.A1(\u_cpu.rf_ram.memory[74][4] ),
    .A2(_02864_),
    .ZN(_02869_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06638_ (.A1(_02748_),
    .A2(_02864_),
    .B(_02869_),
    .ZN(_00251_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06639_ (.A1(\u_cpu.rf_ram.memory[74][5] ),
    .A2(_02864_),
    .ZN(_02870_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06640_ (.A1(_02750_),
    .A2(_02864_),
    .B(_02870_),
    .ZN(_00252_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06641_ (.A1(\u_cpu.rf_ram.memory[74][6] ),
    .A2(_02864_),
    .ZN(_02871_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06642_ (.A1(_02752_),
    .A2(_02864_),
    .B(_02871_),
    .ZN(_00253_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06643_ (.A1(\u_cpu.rf_ram.memory[74][7] ),
    .A2(_02864_),
    .ZN(_02872_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06644_ (.A1(_02754_),
    .A2(_02864_),
    .B(_02872_),
    .ZN(_00254_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06645_ (.A1(_02626_),
    .A2(_02671_),
    .ZN(_02873_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06646_ (.I(_02873_),
    .Z(_02874_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06647_ (.A1(\u_cpu.rf_ram.memory[76][0] ),
    .A2(_02874_),
    .ZN(_02875_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06648_ (.A1(_02738_),
    .A2(_02874_),
    .B(_02875_),
    .ZN(_00255_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06649_ (.A1(\u_cpu.rf_ram.memory[76][1] ),
    .A2(_02874_),
    .ZN(_02876_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06650_ (.A1(_02742_),
    .A2(_02874_),
    .B(_02876_),
    .ZN(_00256_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06651_ (.A1(\u_cpu.rf_ram.memory[76][2] ),
    .A2(_02874_),
    .ZN(_02877_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06652_ (.A1(_02744_),
    .A2(_02874_),
    .B(_02877_),
    .ZN(_00257_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06653_ (.A1(\u_cpu.rf_ram.memory[76][3] ),
    .A2(_02874_),
    .ZN(_02878_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06654_ (.A1(_02746_),
    .A2(_02874_),
    .B(_02878_),
    .ZN(_00258_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06655_ (.A1(\u_cpu.rf_ram.memory[76][4] ),
    .A2(_02874_),
    .ZN(_02879_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06656_ (.A1(_02748_),
    .A2(_02874_),
    .B(_02879_),
    .ZN(_00259_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06657_ (.A1(\u_cpu.rf_ram.memory[76][5] ),
    .A2(_02874_),
    .ZN(_02880_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06658_ (.A1(_02750_),
    .A2(_02874_),
    .B(_02880_),
    .ZN(_00260_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06659_ (.A1(\u_cpu.rf_ram.memory[76][6] ),
    .A2(_02874_),
    .ZN(_02881_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06660_ (.A1(_02752_),
    .A2(_02874_),
    .B(_02881_),
    .ZN(_00261_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06661_ (.A1(\u_cpu.rf_ram.memory[76][7] ),
    .A2(_02874_),
    .ZN(_02882_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06662_ (.A1(_02754_),
    .A2(_02874_),
    .B(_02882_),
    .ZN(_00262_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06663_ (.A1(_02626_),
    .A2(_02706_),
    .ZN(_02883_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06664_ (.I(_02883_),
    .Z(_02884_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06665_ (.A1(\u_cpu.rf_ram.memory[75][0] ),
    .A2(_02884_),
    .ZN(_02885_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06666_ (.A1(_02738_),
    .A2(_02884_),
    .B(_02885_),
    .ZN(_00263_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06667_ (.A1(\u_cpu.rf_ram.memory[75][1] ),
    .A2(_02884_),
    .ZN(_02886_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06668_ (.A1(_02742_),
    .A2(_02884_),
    .B(_02886_),
    .ZN(_00264_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06669_ (.A1(\u_cpu.rf_ram.memory[75][2] ),
    .A2(_02884_),
    .ZN(_02887_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06670_ (.A1(_02744_),
    .A2(_02884_),
    .B(_02887_),
    .ZN(_00265_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06671_ (.A1(\u_cpu.rf_ram.memory[75][3] ),
    .A2(_02884_),
    .ZN(_02888_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06672_ (.A1(_02746_),
    .A2(_02884_),
    .B(_02888_),
    .ZN(_00266_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06673_ (.A1(\u_cpu.rf_ram.memory[75][4] ),
    .A2(_02884_),
    .ZN(_02889_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06674_ (.A1(_02748_),
    .A2(_02884_),
    .B(_02889_),
    .ZN(_00267_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06675_ (.A1(\u_cpu.rf_ram.memory[75][5] ),
    .A2(_02884_),
    .ZN(_02890_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06676_ (.A1(_02750_),
    .A2(_02884_),
    .B(_02890_),
    .ZN(_00268_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06677_ (.A1(\u_cpu.rf_ram.memory[75][6] ),
    .A2(_02884_),
    .ZN(_02891_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06678_ (.A1(_02752_),
    .A2(_02884_),
    .B(_02891_),
    .ZN(_00269_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06679_ (.A1(\u_cpu.rf_ram.memory[75][7] ),
    .A2(_02884_),
    .ZN(_02892_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06680_ (.A1(_02754_),
    .A2(_02884_),
    .B(_02892_),
    .ZN(_00270_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06681_ (.A1(_02468_),
    .A2(_02523_),
    .ZN(_02893_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06682_ (.A1(_02577_),
    .A2(_02893_),
    .ZN(_02894_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06683_ (.I0(_02573_),
    .I1(\u_cpu.rf_ram.memory[6][0] ),
    .S(_02894_),
    .Z(_02895_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06684_ (.I(_02895_),
    .Z(_00271_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06685_ (.I0(_02581_),
    .I1(\u_cpu.rf_ram.memory[6][1] ),
    .S(_02894_),
    .Z(_02896_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06686_ (.I(_02896_),
    .Z(_00272_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06687_ (.I0(_02584_),
    .I1(\u_cpu.rf_ram.memory[6][2] ),
    .S(_02894_),
    .Z(_02897_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06688_ (.I(_02897_),
    .Z(_00273_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06689_ (.I0(_02587_),
    .I1(\u_cpu.rf_ram.memory[6][3] ),
    .S(_02894_),
    .Z(_02898_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06690_ (.I(_02898_),
    .Z(_00274_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06691_ (.I0(_02590_),
    .I1(\u_cpu.rf_ram.memory[6][4] ),
    .S(_02894_),
    .Z(_02899_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06692_ (.I(_02899_),
    .Z(_00275_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06693_ (.I0(_02593_),
    .I1(\u_cpu.rf_ram.memory[6][5] ),
    .S(_02894_),
    .Z(_02900_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06694_ (.I(_02900_),
    .Z(_00276_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06695_ (.I0(_02596_),
    .I1(\u_cpu.rf_ram.memory[6][6] ),
    .S(_02894_),
    .Z(_02901_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06696_ (.I(_02901_),
    .Z(_00277_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06697_ (.I0(_02599_),
    .I1(\u_cpu.rf_ram.memory[6][7] ),
    .S(_02894_),
    .Z(_02902_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06698_ (.I(_02902_),
    .Z(_00278_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06699_ (.A1(_02561_),
    .A2(_02626_),
    .ZN(_02903_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06700_ (.I(_02903_),
    .Z(_02904_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06701_ (.A1(\u_cpu.rf_ram.memory[68][0] ),
    .A2(_02904_),
    .ZN(_02905_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06702_ (.A1(_02738_),
    .A2(_02904_),
    .B(_02905_),
    .ZN(_00279_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06703_ (.A1(\u_cpu.rf_ram.memory[68][1] ),
    .A2(_02904_),
    .ZN(_02906_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06704_ (.A1(_02742_),
    .A2(_02904_),
    .B(_02906_),
    .ZN(_00280_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06705_ (.A1(\u_cpu.rf_ram.memory[68][2] ),
    .A2(_02904_),
    .ZN(_02907_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06706_ (.A1(_02744_),
    .A2(_02904_),
    .B(_02907_),
    .ZN(_00281_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06707_ (.A1(\u_cpu.rf_ram.memory[68][3] ),
    .A2(_02904_),
    .ZN(_02908_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06708_ (.A1(_02746_),
    .A2(_02904_),
    .B(_02908_),
    .ZN(_00282_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06709_ (.A1(\u_cpu.rf_ram.memory[68][4] ),
    .A2(_02904_),
    .ZN(_02909_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06710_ (.A1(_02748_),
    .A2(_02904_),
    .B(_02909_),
    .ZN(_00283_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06711_ (.A1(\u_cpu.rf_ram.memory[68][5] ),
    .A2(_02904_),
    .ZN(_02910_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06712_ (.A1(_02750_),
    .A2(_02904_),
    .B(_02910_),
    .ZN(_00284_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06713_ (.A1(\u_cpu.rf_ram.memory[68][6] ),
    .A2(_02904_),
    .ZN(_02911_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06714_ (.A1(_02752_),
    .A2(_02904_),
    .B(_02911_),
    .ZN(_00285_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06715_ (.A1(\u_cpu.rf_ram.memory[68][7] ),
    .A2(_02904_),
    .ZN(_02912_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06716_ (.A1(_02754_),
    .A2(_02904_),
    .B(_02912_),
    .ZN(_00286_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06717_ (.A1(_02626_),
    .A2(_02682_),
    .ZN(_02913_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06718_ (.I(_02913_),
    .Z(_02914_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06719_ (.A1(\u_cpu.rf_ram.memory[67][0] ),
    .A2(_02914_),
    .ZN(_02915_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06720_ (.A1(_02738_),
    .A2(_02914_),
    .B(_02915_),
    .ZN(_00287_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06721_ (.A1(\u_cpu.rf_ram.memory[67][1] ),
    .A2(_02914_),
    .ZN(_02916_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06722_ (.A1(_02742_),
    .A2(_02914_),
    .B(_02916_),
    .ZN(_00288_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06723_ (.A1(\u_cpu.rf_ram.memory[67][2] ),
    .A2(_02914_),
    .ZN(_02917_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06724_ (.A1(_02744_),
    .A2(_02914_),
    .B(_02917_),
    .ZN(_00289_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06725_ (.A1(\u_cpu.rf_ram.memory[67][3] ),
    .A2(_02914_),
    .ZN(_02918_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06726_ (.A1(_02746_),
    .A2(_02914_),
    .B(_02918_),
    .ZN(_00290_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06727_ (.A1(\u_cpu.rf_ram.memory[67][4] ),
    .A2(_02914_),
    .ZN(_02919_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06728_ (.A1(_02748_),
    .A2(_02914_),
    .B(_02919_),
    .ZN(_00291_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06729_ (.A1(\u_cpu.rf_ram.memory[67][5] ),
    .A2(_02914_),
    .ZN(_02920_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06730_ (.A1(_02750_),
    .A2(_02914_),
    .B(_02920_),
    .ZN(_00292_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06731_ (.A1(\u_cpu.rf_ram.memory[67][6] ),
    .A2(_02914_),
    .ZN(_02921_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06732_ (.A1(_02752_),
    .A2(_02914_),
    .B(_02921_),
    .ZN(_00293_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06733_ (.A1(\u_cpu.rf_ram.memory[67][7] ),
    .A2(_02914_),
    .ZN(_02922_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06734_ (.A1(_02754_),
    .A2(_02914_),
    .B(_02922_),
    .ZN(_00294_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06735_ (.A1(_02469_),
    .A2(_02626_),
    .ZN(_02923_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06736_ (.I(_02923_),
    .Z(_02924_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06737_ (.A1(\u_cpu.rf_ram.memory[66][0] ),
    .A2(_02924_),
    .ZN(_02925_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06738_ (.A1(_02738_),
    .A2(_02924_),
    .B(_02925_),
    .ZN(_00295_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06739_ (.A1(\u_cpu.rf_ram.memory[66][1] ),
    .A2(_02924_),
    .ZN(_02926_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06740_ (.A1(_02742_),
    .A2(_02924_),
    .B(_02926_),
    .ZN(_00296_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06741_ (.A1(\u_cpu.rf_ram.memory[66][2] ),
    .A2(_02924_),
    .ZN(_02927_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06742_ (.A1(_02744_),
    .A2(_02924_),
    .B(_02927_),
    .ZN(_00297_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06743_ (.A1(\u_cpu.rf_ram.memory[66][3] ),
    .A2(_02924_),
    .ZN(_02928_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06744_ (.A1(_02746_),
    .A2(_02924_),
    .B(_02928_),
    .ZN(_00298_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06745_ (.A1(\u_cpu.rf_ram.memory[66][4] ),
    .A2(_02924_),
    .ZN(_02929_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06746_ (.A1(_02748_),
    .A2(_02924_),
    .B(_02929_),
    .ZN(_00299_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06747_ (.A1(\u_cpu.rf_ram.memory[66][5] ),
    .A2(_02924_),
    .ZN(_02930_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06748_ (.A1(_02750_),
    .A2(_02924_),
    .B(_02930_),
    .ZN(_00300_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06749_ (.A1(\u_cpu.rf_ram.memory[66][6] ),
    .A2(_02924_),
    .ZN(_02931_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06750_ (.A1(_02752_),
    .A2(_02924_),
    .B(_02931_),
    .ZN(_00301_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06751_ (.A1(\u_cpu.rf_ram.memory[66][7] ),
    .A2(_02924_),
    .ZN(_02932_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06752_ (.A1(_02754_),
    .A2(_02924_),
    .B(_02932_),
    .ZN(_00302_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06753_ (.A1(_02539_),
    .A2(_02626_),
    .ZN(_02933_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06754_ (.I(_02933_),
    .Z(_02934_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06755_ (.A1(\u_cpu.rf_ram.memory[65][0] ),
    .A2(_02934_),
    .ZN(_02935_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06756_ (.A1(_02738_),
    .A2(_02934_),
    .B(_02935_),
    .ZN(_00303_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06757_ (.A1(\u_cpu.rf_ram.memory[65][1] ),
    .A2(_02934_),
    .ZN(_02936_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06758_ (.A1(_02742_),
    .A2(_02934_),
    .B(_02936_),
    .ZN(_00304_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06759_ (.A1(\u_cpu.rf_ram.memory[65][2] ),
    .A2(_02934_),
    .ZN(_02937_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06760_ (.A1(_02744_),
    .A2(_02934_),
    .B(_02937_),
    .ZN(_00305_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06761_ (.A1(\u_cpu.rf_ram.memory[65][3] ),
    .A2(_02934_),
    .ZN(_02938_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06762_ (.A1(_02746_),
    .A2(_02934_),
    .B(_02938_),
    .ZN(_00306_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06763_ (.A1(\u_cpu.rf_ram.memory[65][4] ),
    .A2(_02934_),
    .ZN(_02939_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06764_ (.A1(_02748_),
    .A2(_02934_),
    .B(_02939_),
    .ZN(_00307_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06765_ (.A1(\u_cpu.rf_ram.memory[65][5] ),
    .A2(_02934_),
    .ZN(_02940_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06766_ (.A1(_02750_),
    .A2(_02934_),
    .B(_02940_),
    .ZN(_00308_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06767_ (.A1(\u_cpu.rf_ram.memory[65][6] ),
    .A2(_02934_),
    .ZN(_02941_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06768_ (.A1(_02752_),
    .A2(_02934_),
    .B(_02941_),
    .ZN(_00309_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06769_ (.A1(\u_cpu.rf_ram.memory[65][7] ),
    .A2(_02934_),
    .ZN(_02942_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06770_ (.A1(_02754_),
    .A2(_02934_),
    .B(_02942_),
    .ZN(_00310_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06771_ (.A1(_02612_),
    .A2(_02626_),
    .ZN(_02943_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06772_ (.I(_02943_),
    .Z(_02944_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06773_ (.A1(\u_cpu.rf_ram.memory[64][0] ),
    .A2(_02944_),
    .ZN(_02945_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06774_ (.A1(_02738_),
    .A2(_02944_),
    .B(_02945_),
    .ZN(_00311_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06775_ (.A1(\u_cpu.rf_ram.memory[64][1] ),
    .A2(_02944_),
    .ZN(_02946_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06776_ (.A1(_02742_),
    .A2(_02944_),
    .B(_02946_),
    .ZN(_00312_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06777_ (.A1(\u_cpu.rf_ram.memory[64][2] ),
    .A2(_02944_),
    .ZN(_02947_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06778_ (.A1(_02744_),
    .A2(_02944_),
    .B(_02947_),
    .ZN(_00313_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06779_ (.A1(\u_cpu.rf_ram.memory[64][3] ),
    .A2(_02944_),
    .ZN(_02948_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06780_ (.A1(_02746_),
    .A2(_02944_),
    .B(_02948_),
    .ZN(_00314_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06781_ (.A1(\u_cpu.rf_ram.memory[64][4] ),
    .A2(_02944_),
    .ZN(_02949_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06782_ (.A1(_02748_),
    .A2(_02944_),
    .B(_02949_),
    .ZN(_00315_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06783_ (.A1(\u_cpu.rf_ram.memory[64][5] ),
    .A2(_02944_),
    .ZN(_02950_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06784_ (.A1(_02750_),
    .A2(_02944_),
    .B(_02950_),
    .ZN(_00316_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06785_ (.A1(\u_cpu.rf_ram.memory[64][6] ),
    .A2(_02944_),
    .ZN(_02951_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06786_ (.A1(_02752_),
    .A2(_02944_),
    .B(_02951_),
    .ZN(_00317_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06787_ (.A1(\u_cpu.rf_ram.memory[64][7] ),
    .A2(_02944_),
    .ZN(_02952_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06788_ (.A1(_02754_),
    .A2(_02944_),
    .B(_02952_),
    .ZN(_00318_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06789_ (.I(_02481_),
    .Z(_02953_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06790_ (.A1(_02528_),
    .A2(_02660_),
    .ZN(_02954_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06791_ (.I(_02954_),
    .Z(_02955_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06792_ (.A1(\u_cpu.rf_ram.memory[29][0] ),
    .A2(_02955_),
    .ZN(_02956_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06793_ (.A1(_02953_),
    .A2(_02955_),
    .B(_02956_),
    .ZN(_00319_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06794_ (.I(_02486_),
    .Z(_02957_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06795_ (.A1(\u_cpu.rf_ram.memory[29][1] ),
    .A2(_02955_),
    .ZN(_02958_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06796_ (.A1(_02957_),
    .A2(_02955_),
    .B(_02958_),
    .ZN(_00320_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06797_ (.I(_02491_),
    .Z(_02959_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06798_ (.A1(\u_cpu.rf_ram.memory[29][2] ),
    .A2(_02955_),
    .ZN(_02960_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06799_ (.A1(_02959_),
    .A2(_02955_),
    .B(_02960_),
    .ZN(_00321_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06800_ (.I(_02496_),
    .Z(_02961_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06801_ (.A1(\u_cpu.rf_ram.memory[29][3] ),
    .A2(_02955_),
    .ZN(_02962_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06802_ (.A1(_02961_),
    .A2(_02955_),
    .B(_02962_),
    .ZN(_00322_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06803_ (.I(_02501_),
    .Z(_02963_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06804_ (.A1(\u_cpu.rf_ram.memory[29][4] ),
    .A2(_02955_),
    .ZN(_02964_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06805_ (.A1(_02963_),
    .A2(_02955_),
    .B(_02964_),
    .ZN(_00323_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06806_ (.I(_02506_),
    .Z(_02965_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06807_ (.A1(\u_cpu.rf_ram.memory[29][5] ),
    .A2(_02955_),
    .ZN(_02966_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06808_ (.A1(_02965_),
    .A2(_02955_),
    .B(_02966_),
    .ZN(_00324_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06809_ (.I(_02511_),
    .Z(_02967_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06810_ (.A1(\u_cpu.rf_ram.memory[29][6] ),
    .A2(_02955_),
    .ZN(_02968_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06811_ (.A1(_02967_),
    .A2(_02955_),
    .B(_02968_),
    .ZN(_00325_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06812_ (.I(_02516_),
    .Z(_02969_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06813_ (.A1(\u_cpu.rf_ram.memory[29][7] ),
    .A2(_02955_),
    .ZN(_02970_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06814_ (.A1(_02969_),
    .A2(_02955_),
    .B(_02970_),
    .ZN(_00326_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06815_ (.A1(_02684_),
    .A2(_02727_),
    .ZN(_02971_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06816_ (.I(_02971_),
    .Z(_02972_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06817_ (.A1(\u_cpu.rf_ram.memory[63][0] ),
    .A2(_02972_),
    .ZN(_02973_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06818_ (.A1(_02953_),
    .A2(_02972_),
    .B(_02973_),
    .ZN(_00327_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06819_ (.A1(\u_cpu.rf_ram.memory[63][1] ),
    .A2(_02972_),
    .ZN(_02974_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06820_ (.A1(_02957_),
    .A2(_02972_),
    .B(_02974_),
    .ZN(_00328_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06821_ (.A1(\u_cpu.rf_ram.memory[63][2] ),
    .A2(_02972_),
    .ZN(_02975_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06822_ (.A1(_02959_),
    .A2(_02972_),
    .B(_02975_),
    .ZN(_00329_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06823_ (.A1(\u_cpu.rf_ram.memory[63][3] ),
    .A2(_02972_),
    .ZN(_02976_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06824_ (.A1(_02961_),
    .A2(_02972_),
    .B(_02976_),
    .ZN(_00330_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06825_ (.A1(\u_cpu.rf_ram.memory[63][4] ),
    .A2(_02972_),
    .ZN(_02977_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06826_ (.A1(_02963_),
    .A2(_02972_),
    .B(_02977_),
    .ZN(_00331_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06827_ (.A1(\u_cpu.rf_ram.memory[63][5] ),
    .A2(_02972_),
    .ZN(_02978_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06828_ (.A1(_02965_),
    .A2(_02972_),
    .B(_02978_),
    .ZN(_00332_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06829_ (.A1(\u_cpu.rf_ram.memory[63][6] ),
    .A2(_02972_),
    .ZN(_02979_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06830_ (.A1(_02967_),
    .A2(_02972_),
    .B(_02979_),
    .ZN(_00333_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06831_ (.A1(\u_cpu.rf_ram.memory[63][7] ),
    .A2(_02972_),
    .ZN(_02980_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06832_ (.A1(_02969_),
    .A2(_02972_),
    .B(_02980_),
    .ZN(_00334_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06833_ (.A1(_02625_),
    .A2(_02684_),
    .ZN(_02981_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06834_ (.I(_02981_),
    .Z(_02982_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06835_ (.A1(\u_cpu.rf_ram.memory[62][0] ),
    .A2(_02982_),
    .ZN(_02983_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06836_ (.A1(_02953_),
    .A2(_02982_),
    .B(_02983_),
    .ZN(_00335_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06837_ (.A1(\u_cpu.rf_ram.memory[62][1] ),
    .A2(_02982_),
    .ZN(_02984_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06838_ (.A1(_02957_),
    .A2(_02982_),
    .B(_02984_),
    .ZN(_00336_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06839_ (.A1(\u_cpu.rf_ram.memory[62][2] ),
    .A2(_02982_),
    .ZN(_02985_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06840_ (.A1(_02959_),
    .A2(_02982_),
    .B(_02985_),
    .ZN(_00337_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06841_ (.A1(\u_cpu.rf_ram.memory[62][3] ),
    .A2(_02982_),
    .ZN(_02986_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06842_ (.A1(_02961_),
    .A2(_02982_),
    .B(_02986_),
    .ZN(_00338_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06843_ (.A1(\u_cpu.rf_ram.memory[62][4] ),
    .A2(_02982_),
    .ZN(_02987_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06844_ (.A1(_02963_),
    .A2(_02982_),
    .B(_02987_),
    .ZN(_00339_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06845_ (.A1(\u_cpu.rf_ram.memory[62][5] ),
    .A2(_02982_),
    .ZN(_02988_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06846_ (.A1(_02965_),
    .A2(_02982_),
    .B(_02988_),
    .ZN(_00340_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06847_ (.A1(\u_cpu.rf_ram.memory[62][6] ),
    .A2(_02982_),
    .ZN(_02989_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06848_ (.A1(_02967_),
    .A2(_02982_),
    .B(_02989_),
    .ZN(_00341_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06849_ (.A1(\u_cpu.rf_ram.memory[62][7] ),
    .A2(_02982_),
    .ZN(_02990_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06850_ (.A1(_02969_),
    .A2(_02982_),
    .B(_02990_),
    .ZN(_00342_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06851_ (.A1(_02660_),
    .A2(_02684_),
    .ZN(_02991_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06852_ (.I(_02991_),
    .Z(_02992_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06853_ (.A1(\u_cpu.rf_ram.memory[61][0] ),
    .A2(_02992_),
    .ZN(_02993_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06854_ (.A1(_02953_),
    .A2(_02992_),
    .B(_02993_),
    .ZN(_00343_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06855_ (.A1(\u_cpu.rf_ram.memory[61][1] ),
    .A2(_02992_),
    .ZN(_02994_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06856_ (.A1(_02957_),
    .A2(_02992_),
    .B(_02994_),
    .ZN(_00344_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06857_ (.A1(\u_cpu.rf_ram.memory[61][2] ),
    .A2(_02992_),
    .ZN(_02995_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06858_ (.A1(_02959_),
    .A2(_02992_),
    .B(_02995_),
    .ZN(_00345_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06859_ (.A1(\u_cpu.rf_ram.memory[61][3] ),
    .A2(_02992_),
    .ZN(_02996_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06860_ (.A1(_02961_),
    .A2(_02992_),
    .B(_02996_),
    .ZN(_00346_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06861_ (.A1(\u_cpu.rf_ram.memory[61][4] ),
    .A2(_02992_),
    .ZN(_02997_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06862_ (.A1(_02963_),
    .A2(_02992_),
    .B(_02997_),
    .ZN(_00347_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06863_ (.A1(\u_cpu.rf_ram.memory[61][5] ),
    .A2(_02992_),
    .ZN(_02998_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06864_ (.A1(_02965_),
    .A2(_02992_),
    .B(_02998_),
    .ZN(_00348_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06865_ (.A1(\u_cpu.rf_ram.memory[61][6] ),
    .A2(_02992_),
    .ZN(_02999_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06866_ (.A1(_02967_),
    .A2(_02992_),
    .B(_02999_),
    .ZN(_00349_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06867_ (.A1(\u_cpu.rf_ram.memory[61][7] ),
    .A2(_02992_),
    .ZN(_03000_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06868_ (.A1(_02969_),
    .A2(_02992_),
    .B(_03000_),
    .ZN(_00350_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06869_ (.A1(_02671_),
    .A2(_02684_),
    .ZN(_03001_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06870_ (.I(_03001_),
    .Z(_03002_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06871_ (.A1(\u_cpu.rf_ram.memory[60][0] ),
    .A2(_03002_),
    .ZN(_03003_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06872_ (.A1(_02953_),
    .A2(_03002_),
    .B(_03003_),
    .ZN(_00351_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06873_ (.A1(\u_cpu.rf_ram.memory[60][1] ),
    .A2(_03002_),
    .ZN(_03004_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06874_ (.A1(_02957_),
    .A2(_03002_),
    .B(_03004_),
    .ZN(_00352_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06875_ (.A1(\u_cpu.rf_ram.memory[60][2] ),
    .A2(_03002_),
    .ZN(_03005_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06876_ (.A1(_02959_),
    .A2(_03002_),
    .B(_03005_),
    .ZN(_00353_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06877_ (.A1(\u_cpu.rf_ram.memory[60][3] ),
    .A2(_03002_),
    .ZN(_03006_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06878_ (.A1(_02961_),
    .A2(_03002_),
    .B(_03006_),
    .ZN(_00354_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06879_ (.A1(\u_cpu.rf_ram.memory[60][4] ),
    .A2(_03002_),
    .ZN(_03007_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06880_ (.A1(_02963_),
    .A2(_03002_),
    .B(_03007_),
    .ZN(_00355_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06881_ (.A1(\u_cpu.rf_ram.memory[60][5] ),
    .A2(_03002_),
    .ZN(_03008_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06882_ (.A1(_02965_),
    .A2(_03002_),
    .B(_03008_),
    .ZN(_00356_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06883_ (.A1(\u_cpu.rf_ram.memory[60][6] ),
    .A2(_03002_),
    .ZN(_03009_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06884_ (.A1(_02967_),
    .A2(_03002_),
    .B(_03009_),
    .ZN(_00357_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06885_ (.A1(\u_cpu.rf_ram.memory[60][7] ),
    .A2(_03002_),
    .ZN(_03010_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06886_ (.A1(_02969_),
    .A2(_03002_),
    .B(_03010_),
    .ZN(_00358_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06887_ (.A1(_02528_),
    .A2(_02682_),
    .ZN(_03011_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06888_ (.I(_03011_),
    .Z(_03012_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06889_ (.A1(\u_cpu.rf_ram.memory[19][0] ),
    .A2(_03012_),
    .ZN(_03013_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06890_ (.A1(_02953_),
    .A2(_03012_),
    .B(_03013_),
    .ZN(_00359_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06891_ (.A1(\u_cpu.rf_ram.memory[19][1] ),
    .A2(_03012_),
    .ZN(_03014_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06892_ (.A1(_02957_),
    .A2(_03012_),
    .B(_03014_),
    .ZN(_00360_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06893_ (.A1(\u_cpu.rf_ram.memory[19][2] ),
    .A2(_03012_),
    .ZN(_03015_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06894_ (.A1(_02959_),
    .A2(_03012_),
    .B(_03015_),
    .ZN(_00361_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06895_ (.A1(\u_cpu.rf_ram.memory[19][3] ),
    .A2(_03012_),
    .ZN(_03016_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06896_ (.A1(_02961_),
    .A2(_03012_),
    .B(_03016_),
    .ZN(_00362_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06897_ (.A1(\u_cpu.rf_ram.memory[19][4] ),
    .A2(_03012_),
    .ZN(_03017_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06898_ (.A1(_02963_),
    .A2(_03012_),
    .B(_03017_),
    .ZN(_00363_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06899_ (.A1(\u_cpu.rf_ram.memory[19][5] ),
    .A2(_03012_),
    .ZN(_03018_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06900_ (.A1(_02965_),
    .A2(_03012_),
    .B(_03018_),
    .ZN(_00364_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06901_ (.A1(\u_cpu.rf_ram.memory[19][6] ),
    .A2(_03012_),
    .ZN(_03019_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06902_ (.A1(_02967_),
    .A2(_03012_),
    .B(_03019_),
    .ZN(_00365_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06903_ (.A1(\u_cpu.rf_ram.memory[19][7] ),
    .A2(_03012_),
    .ZN(_03020_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06904_ (.A1(_02969_),
    .A2(_03012_),
    .B(_03020_),
    .ZN(_00366_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06905_ (.A1(_02524_),
    .A2(_02577_),
    .ZN(_03021_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06906_ (.I0(_02573_),
    .I1(\u_cpu.rf_ram.memory[5][0] ),
    .S(_03021_),
    .Z(_03022_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06907_ (.I(_03022_),
    .Z(_00367_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06908_ (.I0(_02581_),
    .I1(\u_cpu.rf_ram.memory[5][1] ),
    .S(_03021_),
    .Z(_03023_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06909_ (.I(_03023_),
    .Z(_00368_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06910_ (.I0(_02584_),
    .I1(\u_cpu.rf_ram.memory[5][2] ),
    .S(_03021_),
    .Z(_03024_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06911_ (.I(_03024_),
    .Z(_00369_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06912_ (.I0(_02587_),
    .I1(\u_cpu.rf_ram.memory[5][3] ),
    .S(_03021_),
    .Z(_03025_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06913_ (.I(_03025_),
    .Z(_00370_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06914_ (.I0(_02590_),
    .I1(\u_cpu.rf_ram.memory[5][4] ),
    .S(_03021_),
    .Z(_03026_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06915_ (.I(_03026_),
    .Z(_00371_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06916_ (.I0(_02593_),
    .I1(\u_cpu.rf_ram.memory[5][5] ),
    .S(_03021_),
    .Z(_03027_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06917_ (.I(_03027_),
    .Z(_00372_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06918_ (.I0(_02596_),
    .I1(\u_cpu.rf_ram.memory[5][6] ),
    .S(_03021_),
    .Z(_03028_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06919_ (.I(_03028_),
    .Z(_00373_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06920_ (.I0(_02599_),
    .I1(\u_cpu.rf_ram.memory[5][7] ),
    .S(_03021_),
    .Z(_03029_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06921_ (.I(_03029_),
    .Z(_00374_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06922_ (.A1(_02638_),
    .A2(_02684_),
    .ZN(_03030_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06923_ (.I(_03030_),
    .Z(_03031_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06924_ (.A1(\u_cpu.rf_ram.memory[58][0] ),
    .A2(_03031_),
    .ZN(_03032_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06925_ (.A1(_02953_),
    .A2(_03031_),
    .B(_03032_),
    .ZN(_00375_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06926_ (.A1(\u_cpu.rf_ram.memory[58][1] ),
    .A2(_03031_),
    .ZN(_03033_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06927_ (.A1(_02957_),
    .A2(_03031_),
    .B(_03033_),
    .ZN(_00376_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06928_ (.A1(\u_cpu.rf_ram.memory[58][2] ),
    .A2(_03031_),
    .ZN(_03034_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06929_ (.A1(_02959_),
    .A2(_03031_),
    .B(_03034_),
    .ZN(_00377_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06930_ (.A1(\u_cpu.rf_ram.memory[58][3] ),
    .A2(_03031_),
    .ZN(_03035_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06931_ (.A1(_02961_),
    .A2(_03031_),
    .B(_03035_),
    .ZN(_00378_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06932_ (.A1(\u_cpu.rf_ram.memory[58][4] ),
    .A2(_03031_),
    .ZN(_03036_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06933_ (.A1(_02963_),
    .A2(_03031_),
    .B(_03036_),
    .ZN(_00379_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06934_ (.A1(\u_cpu.rf_ram.memory[58][5] ),
    .A2(_03031_),
    .ZN(_03037_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06935_ (.A1(_02965_),
    .A2(_03031_),
    .B(_03037_),
    .ZN(_00380_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06936_ (.A1(\u_cpu.rf_ram.memory[58][6] ),
    .A2(_03031_),
    .ZN(_03038_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06937_ (.A1(_02967_),
    .A2(_03031_),
    .B(_03038_),
    .ZN(_00381_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06938_ (.A1(\u_cpu.rf_ram.memory[58][7] ),
    .A2(_03031_),
    .ZN(_03039_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06939_ (.A1(_02969_),
    .A2(_03031_),
    .B(_03039_),
    .ZN(_00382_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06940_ (.A1(_02684_),
    .A2(_02695_),
    .ZN(_03040_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06941_ (.I(_03040_),
    .Z(_03041_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06942_ (.A1(\u_cpu.rf_ram.memory[57][0] ),
    .A2(_03041_),
    .ZN(_03042_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06943_ (.A1(_02953_),
    .A2(_03041_),
    .B(_03042_),
    .ZN(_00383_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06944_ (.A1(\u_cpu.rf_ram.memory[57][1] ),
    .A2(_03041_),
    .ZN(_03043_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06945_ (.A1(_02957_),
    .A2(_03041_),
    .B(_03043_),
    .ZN(_00384_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06946_ (.A1(\u_cpu.rf_ram.memory[57][2] ),
    .A2(_03041_),
    .ZN(_03044_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06947_ (.A1(_02959_),
    .A2(_03041_),
    .B(_03044_),
    .ZN(_00385_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06948_ (.A1(\u_cpu.rf_ram.memory[57][3] ),
    .A2(_03041_),
    .ZN(_03045_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06949_ (.A1(_02961_),
    .A2(_03041_),
    .B(_03045_),
    .ZN(_00386_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06950_ (.A1(\u_cpu.rf_ram.memory[57][4] ),
    .A2(_03041_),
    .ZN(_03046_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06951_ (.A1(_02963_),
    .A2(_03041_),
    .B(_03046_),
    .ZN(_00387_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06952_ (.A1(\u_cpu.rf_ram.memory[57][5] ),
    .A2(_03041_),
    .ZN(_03047_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06953_ (.A1(_02965_),
    .A2(_03041_),
    .B(_03047_),
    .ZN(_00388_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06954_ (.A1(\u_cpu.rf_ram.memory[57][6] ),
    .A2(_03041_),
    .ZN(_03048_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06955_ (.A1(_02967_),
    .A2(_03041_),
    .B(_03048_),
    .ZN(_00389_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06956_ (.A1(\u_cpu.rf_ram.memory[57][7] ),
    .A2(_03041_),
    .ZN(_03049_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06957_ (.A1(_02969_),
    .A2(_03041_),
    .B(_03049_),
    .ZN(_00390_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06958_ (.A1(_02684_),
    .A2(_02810_),
    .ZN(_03050_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06959_ (.I(_03050_),
    .Z(_03051_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06960_ (.A1(\u_cpu.rf_ram.memory[56][0] ),
    .A2(_03051_),
    .ZN(_03052_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06961_ (.A1(_02953_),
    .A2(_03051_),
    .B(_03052_),
    .ZN(_00391_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06962_ (.A1(\u_cpu.rf_ram.memory[56][1] ),
    .A2(_03051_),
    .ZN(_03053_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06963_ (.A1(_02957_),
    .A2(_03051_),
    .B(_03053_),
    .ZN(_00392_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06964_ (.A1(\u_cpu.rf_ram.memory[56][2] ),
    .A2(_03051_),
    .ZN(_03054_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06965_ (.A1(_02959_),
    .A2(_03051_),
    .B(_03054_),
    .ZN(_00393_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06966_ (.A1(\u_cpu.rf_ram.memory[56][3] ),
    .A2(_03051_),
    .ZN(_03055_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06967_ (.A1(_02961_),
    .A2(_03051_),
    .B(_03055_),
    .ZN(_00394_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06968_ (.A1(\u_cpu.rf_ram.memory[56][4] ),
    .A2(_03051_),
    .ZN(_03056_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06969_ (.A1(_02963_),
    .A2(_03051_),
    .B(_03056_),
    .ZN(_00395_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06970_ (.A1(\u_cpu.rf_ram.memory[56][5] ),
    .A2(_03051_),
    .ZN(_03057_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06971_ (.A1(_02965_),
    .A2(_03051_),
    .B(_03057_),
    .ZN(_00396_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06972_ (.A1(\u_cpu.rf_ram.memory[56][6] ),
    .A2(_03051_),
    .ZN(_03058_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06973_ (.A1(_02967_),
    .A2(_03051_),
    .B(_03058_),
    .ZN(_00397_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06974_ (.A1(\u_cpu.rf_ram.memory[56][7] ),
    .A2(_03051_),
    .ZN(_03059_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06975_ (.A1(_02969_),
    .A2(_03051_),
    .B(_03059_),
    .ZN(_00398_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06976_ (.A1(_02602_),
    .A2(_02684_),
    .ZN(_03060_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06977_ (.I(_03060_),
    .Z(_03061_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06978_ (.A1(\u_cpu.rf_ram.memory[55][0] ),
    .A2(_03061_),
    .ZN(_03062_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06979_ (.A1(_02953_),
    .A2(_03061_),
    .B(_03062_),
    .ZN(_00399_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06980_ (.A1(\u_cpu.rf_ram.memory[55][1] ),
    .A2(_03061_),
    .ZN(_03063_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06981_ (.A1(_02957_),
    .A2(_03061_),
    .B(_03063_),
    .ZN(_00400_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06982_ (.A1(\u_cpu.rf_ram.memory[55][2] ),
    .A2(_03061_),
    .ZN(_03064_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06983_ (.A1(_02959_),
    .A2(_03061_),
    .B(_03064_),
    .ZN(_00401_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06984_ (.A1(\u_cpu.rf_ram.memory[55][3] ),
    .A2(_03061_),
    .ZN(_03065_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06985_ (.A1(_02961_),
    .A2(_03061_),
    .B(_03065_),
    .ZN(_00402_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06986_ (.A1(\u_cpu.rf_ram.memory[55][4] ),
    .A2(_03061_),
    .ZN(_03066_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06987_ (.A1(_02963_),
    .A2(_03061_),
    .B(_03066_),
    .ZN(_00403_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06988_ (.A1(\u_cpu.rf_ram.memory[55][5] ),
    .A2(_03061_),
    .ZN(_03067_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06989_ (.A1(_02965_),
    .A2(_03061_),
    .B(_03067_),
    .ZN(_00404_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06990_ (.A1(\u_cpu.rf_ram.memory[55][6] ),
    .A2(_03061_),
    .ZN(_03068_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06991_ (.A1(_02967_),
    .A2(_03061_),
    .B(_03068_),
    .ZN(_00405_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06992_ (.A1(\u_cpu.rf_ram.memory[55][7] ),
    .A2(_03061_),
    .ZN(_03069_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06993_ (.A1(_02969_),
    .A2(_03061_),
    .B(_03069_),
    .ZN(_00406_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06994_ (.A1(_02684_),
    .A2(_02893_),
    .ZN(_03070_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06995_ (.I(_03070_),
    .Z(_03071_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06996_ (.A1(\u_cpu.rf_ram.memory[54][0] ),
    .A2(_03071_),
    .ZN(_03072_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06997_ (.A1(_02953_),
    .A2(_03071_),
    .B(_03072_),
    .ZN(_00407_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06998_ (.A1(\u_cpu.rf_ram.memory[54][1] ),
    .A2(_03071_),
    .ZN(_03073_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06999_ (.A1(_02957_),
    .A2(_03071_),
    .B(_03073_),
    .ZN(_00408_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07000_ (.A1(\u_cpu.rf_ram.memory[54][2] ),
    .A2(_03071_),
    .ZN(_03074_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07001_ (.A1(_02959_),
    .A2(_03071_),
    .B(_03074_),
    .ZN(_00409_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07002_ (.A1(\u_cpu.rf_ram.memory[54][3] ),
    .A2(_03071_),
    .ZN(_03075_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07003_ (.A1(_02961_),
    .A2(_03071_),
    .B(_03075_),
    .ZN(_00410_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07004_ (.A1(\u_cpu.rf_ram.memory[54][4] ),
    .A2(_03071_),
    .ZN(_03076_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07005_ (.A1(_02963_),
    .A2(_03071_),
    .B(_03076_),
    .ZN(_00411_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07006_ (.A1(\u_cpu.rf_ram.memory[54][5] ),
    .A2(_03071_),
    .ZN(_03077_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07007_ (.A1(_02965_),
    .A2(_03071_),
    .B(_03077_),
    .ZN(_00412_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07008_ (.A1(\u_cpu.rf_ram.memory[54][6] ),
    .A2(_03071_),
    .ZN(_03078_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07009_ (.A1(_02967_),
    .A2(_03071_),
    .B(_03078_),
    .ZN(_00413_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07010_ (.A1(\u_cpu.rf_ram.memory[54][7] ),
    .A2(_03071_),
    .ZN(_03079_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07011_ (.A1(_02969_),
    .A2(_03071_),
    .B(_03079_),
    .ZN(_00414_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07012_ (.A1(_02524_),
    .A2(_02684_),
    .ZN(_03080_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07013_ (.I(_03080_),
    .Z(_03081_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07014_ (.A1(\u_cpu.rf_ram.memory[53][0] ),
    .A2(_03081_),
    .ZN(_03082_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07015_ (.A1(_02953_),
    .A2(_03081_),
    .B(_03082_),
    .ZN(_00415_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07016_ (.A1(\u_cpu.rf_ram.memory[53][1] ),
    .A2(_03081_),
    .ZN(_03083_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07017_ (.A1(_02957_),
    .A2(_03081_),
    .B(_03083_),
    .ZN(_00416_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07018_ (.A1(\u_cpu.rf_ram.memory[53][2] ),
    .A2(_03081_),
    .ZN(_03084_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07019_ (.A1(_02959_),
    .A2(_03081_),
    .B(_03084_),
    .ZN(_00417_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07020_ (.A1(\u_cpu.rf_ram.memory[53][3] ),
    .A2(_03081_),
    .ZN(_03085_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07021_ (.A1(_02961_),
    .A2(_03081_),
    .B(_03085_),
    .ZN(_00418_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07022_ (.A1(\u_cpu.rf_ram.memory[53][4] ),
    .A2(_03081_),
    .ZN(_03086_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07023_ (.A1(_02963_),
    .A2(_03081_),
    .B(_03086_),
    .ZN(_00419_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07024_ (.A1(\u_cpu.rf_ram.memory[53][5] ),
    .A2(_03081_),
    .ZN(_03087_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07025_ (.A1(_02965_),
    .A2(_03081_),
    .B(_03087_),
    .ZN(_00420_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07026_ (.A1(\u_cpu.rf_ram.memory[53][6] ),
    .A2(_03081_),
    .ZN(_03088_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07027_ (.A1(_02967_),
    .A2(_03081_),
    .B(_03088_),
    .ZN(_00421_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07028_ (.A1(\u_cpu.rf_ram.memory[53][7] ),
    .A2(_03081_),
    .ZN(_03089_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07029_ (.A1(_02969_),
    .A2(_03081_),
    .B(_03089_),
    .ZN(_00422_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07030_ (.A1(_02561_),
    .A2(_02684_),
    .ZN(_03090_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07031_ (.I(_03090_),
    .Z(_03091_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07032_ (.A1(\u_cpu.rf_ram.memory[52][0] ),
    .A2(_03091_),
    .ZN(_03092_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07033_ (.A1(_02953_),
    .A2(_03091_),
    .B(_03092_),
    .ZN(_00423_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07034_ (.A1(\u_cpu.rf_ram.memory[52][1] ),
    .A2(_03091_),
    .ZN(_03093_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07035_ (.A1(_02957_),
    .A2(_03091_),
    .B(_03093_),
    .ZN(_00424_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07036_ (.A1(\u_cpu.rf_ram.memory[52][2] ),
    .A2(_03091_),
    .ZN(_03094_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07037_ (.A1(_02959_),
    .A2(_03091_),
    .B(_03094_),
    .ZN(_00425_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07038_ (.A1(\u_cpu.rf_ram.memory[52][3] ),
    .A2(_03091_),
    .ZN(_03095_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07039_ (.A1(_02961_),
    .A2(_03091_),
    .B(_03095_),
    .ZN(_00426_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07040_ (.A1(\u_cpu.rf_ram.memory[52][4] ),
    .A2(_03091_),
    .ZN(_03096_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07041_ (.A1(_02963_),
    .A2(_03091_),
    .B(_03096_),
    .ZN(_00427_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07042_ (.A1(\u_cpu.rf_ram.memory[52][5] ),
    .A2(_03091_),
    .ZN(_03097_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07043_ (.A1(_02965_),
    .A2(_03091_),
    .B(_03097_),
    .ZN(_00428_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07044_ (.A1(\u_cpu.rf_ram.memory[52][6] ),
    .A2(_03091_),
    .ZN(_03098_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07045_ (.A1(_02967_),
    .A2(_03091_),
    .B(_03098_),
    .ZN(_00429_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07046_ (.A1(\u_cpu.rf_ram.memory[52][7] ),
    .A2(_03091_),
    .ZN(_03099_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07047_ (.A1(_02969_),
    .A2(_03091_),
    .B(_03099_),
    .ZN(_00430_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07048_ (.A1(_02577_),
    .A2(_02695_),
    .ZN(_03100_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07049_ (.I0(_02573_),
    .I1(\u_cpu.rf_ram.memory[9][0] ),
    .S(_03100_),
    .Z(_03101_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07050_ (.I(_03101_),
    .Z(_00431_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07051_ (.I0(_02581_),
    .I1(\u_cpu.rf_ram.memory[9][1] ),
    .S(_03100_),
    .Z(_03102_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07052_ (.I(_03102_),
    .Z(_00432_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07053_ (.I0(_02584_),
    .I1(\u_cpu.rf_ram.memory[9][2] ),
    .S(_03100_),
    .Z(_03103_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07054_ (.I(_03103_),
    .Z(_00433_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07055_ (.I0(_02587_),
    .I1(\u_cpu.rf_ram.memory[9][3] ),
    .S(_03100_),
    .Z(_03104_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07056_ (.I(_03104_),
    .Z(_00434_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07057_ (.I0(_02590_),
    .I1(\u_cpu.rf_ram.memory[9][4] ),
    .S(_03100_),
    .Z(_03105_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07058_ (.I(_03105_),
    .Z(_00435_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07059_ (.I0(_02593_),
    .I1(\u_cpu.rf_ram.memory[9][5] ),
    .S(_03100_),
    .Z(_03106_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07060_ (.I(_03106_),
    .Z(_00436_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07061_ (.I0(_02596_),
    .I1(\u_cpu.rf_ram.memory[9][6] ),
    .S(_03100_),
    .Z(_03107_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07062_ (.I(_03107_),
    .Z(_00437_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07063_ (.I0(_02599_),
    .I1(\u_cpu.rf_ram.memory[9][7] ),
    .S(_03100_),
    .Z(_03108_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07064_ (.I(_03108_),
    .Z(_00438_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07065_ (.A1(_02577_),
    .A2(_02727_),
    .ZN(_03109_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07066_ (.I0(_02573_),
    .I1(\u_cpu.rf_ram.memory[15][0] ),
    .S(_03109_),
    .Z(_03110_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07067_ (.I(_03110_),
    .Z(_00439_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07068_ (.I0(_02581_),
    .I1(\u_cpu.rf_ram.memory[15][1] ),
    .S(_03109_),
    .Z(_03111_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07069_ (.I(_03111_),
    .Z(_00440_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07070_ (.I0(_02584_),
    .I1(\u_cpu.rf_ram.memory[15][2] ),
    .S(_03109_),
    .Z(_03112_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07071_ (.I(_03112_),
    .Z(_00441_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07072_ (.I0(_02587_),
    .I1(\u_cpu.rf_ram.memory[15][3] ),
    .S(_03109_),
    .Z(_03113_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07073_ (.I(_03113_),
    .Z(_00442_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07074_ (.I0(_02590_),
    .I1(\u_cpu.rf_ram.memory[15][4] ),
    .S(_03109_),
    .Z(_03114_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07075_ (.I(_03114_),
    .Z(_00443_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07076_ (.I0(_02593_),
    .I1(\u_cpu.rf_ram.memory[15][5] ),
    .S(_03109_),
    .Z(_03115_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07077_ (.I(_03115_),
    .Z(_00444_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07078_ (.I0(_02596_),
    .I1(\u_cpu.rf_ram.memory[15][6] ),
    .S(_03109_),
    .Z(_03116_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07079_ (.I(_03116_),
    .Z(_00445_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07080_ (.I0(_02599_),
    .I1(\u_cpu.rf_ram.memory[15][7] ),
    .S(_03109_),
    .Z(_03117_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07081_ (.I(_03117_),
    .Z(_00446_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07082_ (.A1(_02625_),
    .A2(_02832_),
    .ZN(_03118_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07083_ (.I(_03118_),
    .Z(_03119_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07084_ (.A1(\u_cpu.rf_ram.memory[142][0] ),
    .A2(_03119_),
    .ZN(_03120_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07085_ (.A1(_02953_),
    .A2(_03119_),
    .B(_03120_),
    .ZN(_00447_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07086_ (.A1(\u_cpu.rf_ram.memory[142][1] ),
    .A2(_03119_),
    .ZN(_03121_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07087_ (.A1(_02957_),
    .A2(_03119_),
    .B(_03121_),
    .ZN(_00448_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07088_ (.A1(\u_cpu.rf_ram.memory[142][2] ),
    .A2(_03119_),
    .ZN(_03122_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07089_ (.A1(_02959_),
    .A2(_03119_),
    .B(_03122_),
    .ZN(_00449_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07090_ (.A1(\u_cpu.rf_ram.memory[142][3] ),
    .A2(_03119_),
    .ZN(_03123_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07091_ (.A1(_02961_),
    .A2(_03119_),
    .B(_03123_),
    .ZN(_00450_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07092_ (.A1(\u_cpu.rf_ram.memory[142][4] ),
    .A2(_03119_),
    .ZN(_03124_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07093_ (.A1(_02963_),
    .A2(_03119_),
    .B(_03124_),
    .ZN(_00451_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07094_ (.A1(\u_cpu.rf_ram.memory[142][5] ),
    .A2(_03119_),
    .ZN(_03125_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07095_ (.A1(_02965_),
    .A2(_03119_),
    .B(_03125_),
    .ZN(_00452_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07096_ (.A1(\u_cpu.rf_ram.memory[142][6] ),
    .A2(_03119_),
    .ZN(_03126_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07097_ (.A1(_02967_),
    .A2(_03119_),
    .B(_03126_),
    .ZN(_00453_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07098_ (.A1(\u_cpu.rf_ram.memory[142][7] ),
    .A2(_03119_),
    .ZN(_03127_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07099_ (.A1(_02969_),
    .A2(_03119_),
    .B(_03127_),
    .ZN(_00454_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07100_ (.A1(_02660_),
    .A2(_02832_),
    .ZN(_03128_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07101_ (.I(_03128_),
    .Z(_03129_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07102_ (.A1(\u_cpu.rf_ram.memory[141][0] ),
    .A2(_03129_),
    .ZN(_03130_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07103_ (.A1(_02953_),
    .A2(_03129_),
    .B(_03130_),
    .ZN(_00455_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07104_ (.A1(\u_cpu.rf_ram.memory[141][1] ),
    .A2(_03129_),
    .ZN(_03131_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07105_ (.A1(_02957_),
    .A2(_03129_),
    .B(_03131_),
    .ZN(_00456_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07106_ (.A1(\u_cpu.rf_ram.memory[141][2] ),
    .A2(_03129_),
    .ZN(_03132_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07107_ (.A1(_02959_),
    .A2(_03129_),
    .B(_03132_),
    .ZN(_00457_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07108_ (.A1(\u_cpu.rf_ram.memory[141][3] ),
    .A2(_03129_),
    .ZN(_03133_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07109_ (.A1(_02961_),
    .A2(_03129_),
    .B(_03133_),
    .ZN(_00458_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07110_ (.A1(\u_cpu.rf_ram.memory[141][4] ),
    .A2(_03129_),
    .ZN(_03134_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07111_ (.A1(_02963_),
    .A2(_03129_),
    .B(_03134_),
    .ZN(_00459_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07112_ (.A1(\u_cpu.rf_ram.memory[141][5] ),
    .A2(_03129_),
    .ZN(_03135_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07113_ (.A1(_02965_),
    .A2(_03129_),
    .B(_03135_),
    .ZN(_00460_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07114_ (.A1(\u_cpu.rf_ram.memory[141][6] ),
    .A2(_03129_),
    .ZN(_03136_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07115_ (.A1(_02967_),
    .A2(_03129_),
    .B(_03136_),
    .ZN(_00461_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07116_ (.A1(\u_cpu.rf_ram.memory[141][7] ),
    .A2(_03129_),
    .ZN(_03137_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07117_ (.A1(_02969_),
    .A2(_03129_),
    .B(_03137_),
    .ZN(_00462_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07118_ (.A1(_02671_),
    .A2(_02832_),
    .ZN(_03138_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07119_ (.I(_03138_),
    .Z(_03139_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07120_ (.A1(\u_cpu.rf_ram.memory[140][0] ),
    .A2(_03139_),
    .ZN(_03140_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07121_ (.A1(_02953_),
    .A2(_03139_),
    .B(_03140_),
    .ZN(_00463_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07122_ (.A1(\u_cpu.rf_ram.memory[140][1] ),
    .A2(_03139_),
    .ZN(_03141_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07123_ (.A1(_02957_),
    .A2(_03139_),
    .B(_03141_),
    .ZN(_00464_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07124_ (.A1(\u_cpu.rf_ram.memory[140][2] ),
    .A2(_03139_),
    .ZN(_03142_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07125_ (.A1(_02959_),
    .A2(_03139_),
    .B(_03142_),
    .ZN(_00465_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07126_ (.A1(\u_cpu.rf_ram.memory[140][3] ),
    .A2(_03139_),
    .ZN(_03143_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07127_ (.A1(_02961_),
    .A2(_03139_),
    .B(_03143_),
    .ZN(_00466_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07128_ (.A1(\u_cpu.rf_ram.memory[140][4] ),
    .A2(_03139_),
    .ZN(_03144_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07129_ (.A1(_02963_),
    .A2(_03139_),
    .B(_03144_),
    .ZN(_00467_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07130_ (.A1(\u_cpu.rf_ram.memory[140][5] ),
    .A2(_03139_),
    .ZN(_03145_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07131_ (.A1(_02965_),
    .A2(_03139_),
    .B(_03145_),
    .ZN(_00468_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07132_ (.A1(\u_cpu.rf_ram.memory[140][6] ),
    .A2(_03139_),
    .ZN(_03146_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07133_ (.A1(_02967_),
    .A2(_03139_),
    .B(_03146_),
    .ZN(_00469_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07134_ (.A1(\u_cpu.rf_ram.memory[140][7] ),
    .A2(_03139_),
    .ZN(_03147_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07135_ (.A1(_02969_),
    .A2(_03139_),
    .B(_03147_),
    .ZN(_00470_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07136_ (.A1(_02577_),
    .A2(_02660_),
    .ZN(_03148_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07137_ (.I0(_02573_),
    .I1(\u_cpu.rf_ram.memory[13][0] ),
    .S(_03148_),
    .Z(_03149_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07138_ (.I(_03149_),
    .Z(_00471_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07139_ (.I0(_02581_),
    .I1(\u_cpu.rf_ram.memory[13][1] ),
    .S(_03148_),
    .Z(_03150_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07140_ (.I(_03150_),
    .Z(_00472_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07141_ (.I0(_02584_),
    .I1(\u_cpu.rf_ram.memory[13][2] ),
    .S(_03148_),
    .Z(_03151_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07142_ (.I(_03151_),
    .Z(_00473_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07143_ (.I0(_02587_),
    .I1(\u_cpu.rf_ram.memory[13][3] ),
    .S(_03148_),
    .Z(_03152_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07144_ (.I(_03152_),
    .Z(_00474_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07145_ (.I0(_02590_),
    .I1(\u_cpu.rf_ram.memory[13][4] ),
    .S(_03148_),
    .Z(_03153_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07146_ (.I(_03153_),
    .Z(_00475_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07147_ (.I0(_02593_),
    .I1(\u_cpu.rf_ram.memory[13][5] ),
    .S(_03148_),
    .Z(_03154_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07148_ (.I(_03154_),
    .Z(_00476_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07149_ (.I0(_02596_),
    .I1(\u_cpu.rf_ram.memory[13][6] ),
    .S(_03148_),
    .Z(_03155_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07150_ (.I(_03155_),
    .Z(_00477_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07151_ (.I0(_02599_),
    .I1(\u_cpu.rf_ram.memory[13][7] ),
    .S(_03148_),
    .Z(_03156_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07152_ (.I(_03156_),
    .Z(_00478_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07153_ (.I(_02481_),
    .Z(_03157_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07154_ (.A1(_02626_),
    .A2(_02810_),
    .ZN(_03158_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07155_ (.I(_03158_),
    .Z(_03159_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07156_ (.A1(\u_cpu.rf_ram.memory[72][0] ),
    .A2(_03159_),
    .ZN(_03160_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07157_ (.A1(_03157_),
    .A2(_03159_),
    .B(_03160_),
    .ZN(_00479_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07158_ (.I(_02486_),
    .Z(_03161_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07159_ (.A1(\u_cpu.rf_ram.memory[72][1] ),
    .A2(_03159_),
    .ZN(_03162_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07160_ (.A1(_03161_),
    .A2(_03159_),
    .B(_03162_),
    .ZN(_00480_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07161_ (.I(_02491_),
    .Z(_03163_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07162_ (.A1(\u_cpu.rf_ram.memory[72][2] ),
    .A2(_03159_),
    .ZN(_03164_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07163_ (.A1(_03163_),
    .A2(_03159_),
    .B(_03164_),
    .ZN(_00481_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07164_ (.I(_02496_),
    .Z(_03165_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07165_ (.A1(\u_cpu.rf_ram.memory[72][3] ),
    .A2(_03159_),
    .ZN(_03166_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07166_ (.A1(_03165_),
    .A2(_03159_),
    .B(_03166_),
    .ZN(_00482_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07167_ (.I(_02501_),
    .Z(_03167_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07168_ (.A1(\u_cpu.rf_ram.memory[72][4] ),
    .A2(_03159_),
    .ZN(_03168_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07169_ (.A1(_03167_),
    .A2(_03159_),
    .B(_03168_),
    .ZN(_00483_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07170_ (.I(_02506_),
    .Z(_03169_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07171_ (.A1(\u_cpu.rf_ram.memory[72][5] ),
    .A2(_03159_),
    .ZN(_03170_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07172_ (.A1(_03169_),
    .A2(_03159_),
    .B(_03170_),
    .ZN(_00484_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07173_ (.I(_02511_),
    .Z(_03171_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07174_ (.A1(\u_cpu.rf_ram.memory[72][6] ),
    .A2(_03159_),
    .ZN(_03172_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07175_ (.A1(_03171_),
    .A2(_03159_),
    .B(_03172_),
    .ZN(_00485_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07176_ (.I(_02516_),
    .Z(_03173_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07177_ (.A1(\u_cpu.rf_ram.memory[72][7] ),
    .A2(_03159_),
    .ZN(_03174_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07178_ (.A1(_03173_),
    .A2(_03159_),
    .B(_03174_),
    .ZN(_00486_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07179_ (.A1(_02626_),
    .A2(_02695_),
    .ZN(_03175_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07180_ (.I(_03175_),
    .Z(_03176_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07181_ (.A1(\u_cpu.rf_ram.memory[73][0] ),
    .A2(_03176_),
    .ZN(_03177_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07182_ (.A1(_03157_),
    .A2(_03176_),
    .B(_03177_),
    .ZN(_00487_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07183_ (.A1(\u_cpu.rf_ram.memory[73][1] ),
    .A2(_03176_),
    .ZN(_03178_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07184_ (.A1(_03161_),
    .A2(_03176_),
    .B(_03178_),
    .ZN(_00488_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07185_ (.A1(\u_cpu.rf_ram.memory[73][2] ),
    .A2(_03176_),
    .ZN(_03179_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07186_ (.A1(_03163_),
    .A2(_03176_),
    .B(_03179_),
    .ZN(_00489_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07187_ (.A1(\u_cpu.rf_ram.memory[73][3] ),
    .A2(_03176_),
    .ZN(_03180_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07188_ (.A1(_03165_),
    .A2(_03176_),
    .B(_03180_),
    .ZN(_00490_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07189_ (.A1(\u_cpu.rf_ram.memory[73][4] ),
    .A2(_03176_),
    .ZN(_03181_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07190_ (.A1(_03167_),
    .A2(_03176_),
    .B(_03181_),
    .ZN(_00491_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07191_ (.A1(\u_cpu.rf_ram.memory[73][5] ),
    .A2(_03176_),
    .ZN(_03182_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07192_ (.A1(_03169_),
    .A2(_03176_),
    .B(_03182_),
    .ZN(_00492_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07193_ (.A1(\u_cpu.rf_ram.memory[73][6] ),
    .A2(_03176_),
    .ZN(_03183_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07194_ (.A1(_03171_),
    .A2(_03176_),
    .B(_03183_),
    .ZN(_00493_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07195_ (.A1(\u_cpu.rf_ram.memory[73][7] ),
    .A2(_03176_),
    .ZN(_03184_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07196_ (.A1(_03173_),
    .A2(_03176_),
    .B(_03184_),
    .ZN(_00494_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07197_ (.A1(_02602_),
    .A2(_02626_),
    .ZN(_03185_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07198_ (.I(_03185_),
    .Z(_03186_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07199_ (.A1(\u_cpu.rf_ram.memory[71][0] ),
    .A2(_03186_),
    .ZN(_03187_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07200_ (.A1(_03157_),
    .A2(_03186_),
    .B(_03187_),
    .ZN(_00495_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07201_ (.A1(\u_cpu.rf_ram.memory[71][1] ),
    .A2(_03186_),
    .ZN(_03188_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07202_ (.A1(_03161_),
    .A2(_03186_),
    .B(_03188_),
    .ZN(_00496_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07203_ (.A1(\u_cpu.rf_ram.memory[71][2] ),
    .A2(_03186_),
    .ZN(_03189_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07204_ (.A1(_03163_),
    .A2(_03186_),
    .B(_03189_),
    .ZN(_00497_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07205_ (.A1(\u_cpu.rf_ram.memory[71][3] ),
    .A2(_03186_),
    .ZN(_03190_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07206_ (.A1(_03165_),
    .A2(_03186_),
    .B(_03190_),
    .ZN(_00498_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07207_ (.A1(\u_cpu.rf_ram.memory[71][4] ),
    .A2(_03186_),
    .ZN(_03191_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07208_ (.A1(_03167_),
    .A2(_03186_),
    .B(_03191_),
    .ZN(_00499_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07209_ (.A1(\u_cpu.rf_ram.memory[71][5] ),
    .A2(_03186_),
    .ZN(_03192_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07210_ (.A1(_03169_),
    .A2(_03186_),
    .B(_03192_),
    .ZN(_00500_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07211_ (.A1(\u_cpu.rf_ram.memory[71][6] ),
    .A2(_03186_),
    .ZN(_03193_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07212_ (.A1(_03171_),
    .A2(_03186_),
    .B(_03193_),
    .ZN(_00501_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07213_ (.A1(\u_cpu.rf_ram.memory[71][7] ),
    .A2(_03186_),
    .ZN(_03194_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07214_ (.A1(_03173_),
    .A2(_03186_),
    .B(_03194_),
    .ZN(_00502_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07215_ (.A1(_02626_),
    .A2(_02893_),
    .ZN(_03195_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07216_ (.I(_03195_),
    .Z(_03196_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07217_ (.A1(\u_cpu.rf_ram.memory[70][0] ),
    .A2(_03196_),
    .ZN(_03197_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07218_ (.A1(_03157_),
    .A2(_03196_),
    .B(_03197_),
    .ZN(_00503_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07219_ (.A1(\u_cpu.rf_ram.memory[70][1] ),
    .A2(_03196_),
    .ZN(_03198_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07220_ (.A1(_03161_),
    .A2(_03196_),
    .B(_03198_),
    .ZN(_00504_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07221_ (.A1(\u_cpu.rf_ram.memory[70][2] ),
    .A2(_03196_),
    .ZN(_03199_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07222_ (.A1(_03163_),
    .A2(_03196_),
    .B(_03199_),
    .ZN(_00505_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07223_ (.A1(\u_cpu.rf_ram.memory[70][3] ),
    .A2(_03196_),
    .ZN(_03200_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07224_ (.A1(_03165_),
    .A2(_03196_),
    .B(_03200_),
    .ZN(_00506_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07225_ (.A1(\u_cpu.rf_ram.memory[70][4] ),
    .A2(_03196_),
    .ZN(_03201_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07226_ (.A1(_03167_),
    .A2(_03196_),
    .B(_03201_),
    .ZN(_00507_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07227_ (.A1(\u_cpu.rf_ram.memory[70][5] ),
    .A2(_03196_),
    .ZN(_03202_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07228_ (.A1(_03169_),
    .A2(_03196_),
    .B(_03202_),
    .ZN(_00508_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07229_ (.A1(\u_cpu.rf_ram.memory[70][6] ),
    .A2(_03196_),
    .ZN(_03203_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07230_ (.A1(_03171_),
    .A2(_03196_),
    .B(_03203_),
    .ZN(_00509_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07231_ (.A1(\u_cpu.rf_ram.memory[70][7] ),
    .A2(_03196_),
    .ZN(_03204_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07232_ (.A1(_03173_),
    .A2(_03196_),
    .B(_03204_),
    .ZN(_00510_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07233_ (.A1(_02727_),
    .A2(_02832_),
    .ZN(_03205_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07234_ (.I(_03205_),
    .Z(_03206_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07235_ (.A1(\u_cpu.rf_ram.memory[143][0] ),
    .A2(_03206_),
    .ZN(_03207_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07236_ (.A1(_03157_),
    .A2(_03206_),
    .B(_03207_),
    .ZN(_00511_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07237_ (.A1(\u_cpu.rf_ram.memory[143][1] ),
    .A2(_03206_),
    .ZN(_03208_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07238_ (.A1(_03161_),
    .A2(_03206_),
    .B(_03208_),
    .ZN(_00512_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07239_ (.A1(\u_cpu.rf_ram.memory[143][2] ),
    .A2(_03206_),
    .ZN(_03209_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07240_ (.A1(_03163_),
    .A2(_03206_),
    .B(_03209_),
    .ZN(_00513_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07241_ (.A1(\u_cpu.rf_ram.memory[143][3] ),
    .A2(_03206_),
    .ZN(_03210_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07242_ (.A1(_03165_),
    .A2(_03206_),
    .B(_03210_),
    .ZN(_00514_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07243_ (.A1(\u_cpu.rf_ram.memory[143][4] ),
    .A2(_03206_),
    .ZN(_03211_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07244_ (.A1(_03167_),
    .A2(_03206_),
    .B(_03211_),
    .ZN(_00515_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07245_ (.A1(\u_cpu.rf_ram.memory[143][5] ),
    .A2(_03206_),
    .ZN(_03212_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07246_ (.A1(_03169_),
    .A2(_03206_),
    .B(_03212_),
    .ZN(_00516_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07247_ (.A1(\u_cpu.rf_ram.memory[143][6] ),
    .A2(_03206_),
    .ZN(_03213_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07248_ (.A1(_03171_),
    .A2(_03206_),
    .B(_03213_),
    .ZN(_00517_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07249_ (.A1(\u_cpu.rf_ram.memory[143][7] ),
    .A2(_03206_),
    .ZN(_03214_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07250_ (.A1(_03173_),
    .A2(_03206_),
    .B(_03214_),
    .ZN(_00518_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07251_ (.A1(_02577_),
    .A2(_02625_),
    .ZN(_03215_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07252_ (.I0(_02573_),
    .I1(\u_cpu.rf_ram.memory[14][0] ),
    .S(_03215_),
    .Z(_03216_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07253_ (.I(_03216_),
    .Z(_00519_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07254_ (.I0(_02581_),
    .I1(\u_cpu.rf_ram.memory[14][1] ),
    .S(_03215_),
    .Z(_03217_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07255_ (.I(_03217_),
    .Z(_00520_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07256_ (.I0(_02584_),
    .I1(\u_cpu.rf_ram.memory[14][2] ),
    .S(_03215_),
    .Z(_03218_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07257_ (.I(_03218_),
    .Z(_00521_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07258_ (.I0(_02587_),
    .I1(\u_cpu.rf_ram.memory[14][3] ),
    .S(_03215_),
    .Z(_03219_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07259_ (.I(_03219_),
    .Z(_00522_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07260_ (.I0(_02590_),
    .I1(\u_cpu.rf_ram.memory[14][4] ),
    .S(_03215_),
    .Z(_03220_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07261_ (.I(_03220_),
    .Z(_00523_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07262_ (.I0(_02593_),
    .I1(\u_cpu.rf_ram.memory[14][5] ),
    .S(_03215_),
    .Z(_03221_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07263_ (.I(_03221_),
    .Z(_00524_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07264_ (.I0(_02596_),
    .I1(\u_cpu.rf_ram.memory[14][6] ),
    .S(_03215_),
    .Z(_03222_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07265_ (.I(_03222_),
    .Z(_00525_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07266_ (.I0(_02599_),
    .I1(\u_cpu.rf_ram.memory[14][7] ),
    .S(_03215_),
    .Z(_03223_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07267_ (.I(_03223_),
    .Z(_00526_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07268_ (.A1(_02638_),
    .A2(_02832_),
    .ZN(_03224_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07269_ (.I(_03224_),
    .Z(_03225_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07270_ (.A1(\u_cpu.rf_ram.memory[138][0] ),
    .A2(_03225_),
    .ZN(_03226_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07271_ (.A1(_03157_),
    .A2(_03225_),
    .B(_03226_),
    .ZN(_00527_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07272_ (.A1(\u_cpu.rf_ram.memory[138][1] ),
    .A2(_03225_),
    .ZN(_03227_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07273_ (.A1(_03161_),
    .A2(_03225_),
    .B(_03227_),
    .ZN(_00528_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07274_ (.A1(\u_cpu.rf_ram.memory[138][2] ),
    .A2(_03225_),
    .ZN(_03228_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07275_ (.A1(_03163_),
    .A2(_03225_),
    .B(_03228_),
    .ZN(_00529_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07276_ (.A1(\u_cpu.rf_ram.memory[138][3] ),
    .A2(_03225_),
    .ZN(_03229_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07277_ (.A1(_03165_),
    .A2(_03225_),
    .B(_03229_),
    .ZN(_00530_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07278_ (.A1(\u_cpu.rf_ram.memory[138][4] ),
    .A2(_03225_),
    .ZN(_03230_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07279_ (.A1(_03167_),
    .A2(_03225_),
    .B(_03230_),
    .ZN(_00531_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07280_ (.A1(\u_cpu.rf_ram.memory[138][5] ),
    .A2(_03225_),
    .ZN(_03231_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07281_ (.A1(_03169_),
    .A2(_03225_),
    .B(_03231_),
    .ZN(_00532_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07282_ (.A1(\u_cpu.rf_ram.memory[138][6] ),
    .A2(_03225_),
    .ZN(_03232_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07283_ (.A1(_03171_),
    .A2(_03225_),
    .B(_03232_),
    .ZN(_00533_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07284_ (.A1(\u_cpu.rf_ram.memory[138][7] ),
    .A2(_03225_),
    .ZN(_03233_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07285_ (.A1(_03173_),
    .A2(_03225_),
    .B(_03233_),
    .ZN(_00534_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07286_ (.A1(_02602_),
    .A2(_02639_),
    .ZN(_03234_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07287_ (.I(_03234_),
    .Z(_03235_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07288_ (.A1(\u_cpu.rf_ram.memory[39][0] ),
    .A2(_03235_),
    .ZN(_03236_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07289_ (.A1(_03157_),
    .A2(_03235_),
    .B(_03236_),
    .ZN(_00535_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07290_ (.A1(\u_cpu.rf_ram.memory[39][1] ),
    .A2(_03235_),
    .ZN(_03237_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07291_ (.A1(_03161_),
    .A2(_03235_),
    .B(_03237_),
    .ZN(_00536_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07292_ (.A1(\u_cpu.rf_ram.memory[39][2] ),
    .A2(_03235_),
    .ZN(_03238_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07293_ (.A1(_03163_),
    .A2(_03235_),
    .B(_03238_),
    .ZN(_00537_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07294_ (.A1(\u_cpu.rf_ram.memory[39][3] ),
    .A2(_03235_),
    .ZN(_03239_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07295_ (.A1(_03165_),
    .A2(_03235_),
    .B(_03239_),
    .ZN(_00538_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07296_ (.A1(\u_cpu.rf_ram.memory[39][4] ),
    .A2(_03235_),
    .ZN(_03240_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07297_ (.A1(_03167_),
    .A2(_03235_),
    .B(_03240_),
    .ZN(_00539_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07298_ (.A1(\u_cpu.rf_ram.memory[39][5] ),
    .A2(_03235_),
    .ZN(_03241_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07299_ (.A1(_03169_),
    .A2(_03235_),
    .B(_03241_),
    .ZN(_00540_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07300_ (.A1(\u_cpu.rf_ram.memory[39][6] ),
    .A2(_03235_),
    .ZN(_03242_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07301_ (.A1(_03171_),
    .A2(_03235_),
    .B(_03242_),
    .ZN(_00541_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07302_ (.A1(\u_cpu.rf_ram.memory[39][7] ),
    .A2(_03235_),
    .ZN(_03243_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07303_ (.A1(_03173_),
    .A2(_03235_),
    .B(_03243_),
    .ZN(_00542_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07304_ (.A1(_02695_),
    .A2(_02832_),
    .ZN(_03244_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07305_ (.I(_03244_),
    .Z(_03245_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07306_ (.A1(\u_cpu.rf_ram.memory[137][0] ),
    .A2(_03245_),
    .ZN(_03246_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07307_ (.A1(_03157_),
    .A2(_03245_),
    .B(_03246_),
    .ZN(_00543_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07308_ (.A1(\u_cpu.rf_ram.memory[137][1] ),
    .A2(_03245_),
    .ZN(_03247_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07309_ (.A1(_03161_),
    .A2(_03245_),
    .B(_03247_),
    .ZN(_00544_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07310_ (.A1(\u_cpu.rf_ram.memory[137][2] ),
    .A2(_03245_),
    .ZN(_03248_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07311_ (.A1(_03163_),
    .A2(_03245_),
    .B(_03248_),
    .ZN(_00545_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07312_ (.A1(\u_cpu.rf_ram.memory[137][3] ),
    .A2(_03245_),
    .ZN(_03249_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07313_ (.A1(_03165_),
    .A2(_03245_),
    .B(_03249_),
    .ZN(_00546_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07314_ (.A1(\u_cpu.rf_ram.memory[137][4] ),
    .A2(_03245_),
    .ZN(_03250_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07315_ (.A1(_03167_),
    .A2(_03245_),
    .B(_03250_),
    .ZN(_00547_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07316_ (.A1(\u_cpu.rf_ram.memory[137][5] ),
    .A2(_03245_),
    .ZN(_03251_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07317_ (.A1(_03169_),
    .A2(_03245_),
    .B(_03251_),
    .ZN(_00548_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07318_ (.A1(\u_cpu.rf_ram.memory[137][6] ),
    .A2(_03245_),
    .ZN(_03252_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07319_ (.A1(_03171_),
    .A2(_03245_),
    .B(_03252_),
    .ZN(_00549_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07320_ (.A1(\u_cpu.rf_ram.memory[137][7] ),
    .A2(_03245_),
    .ZN(_03253_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07321_ (.A1(_03173_),
    .A2(_03245_),
    .B(_03253_),
    .ZN(_00550_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07322_ (.A1(_02539_),
    .A2(_02684_),
    .ZN(_03254_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07323_ (.I(_03254_),
    .Z(_03255_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07324_ (.A1(\u_cpu.rf_ram.memory[49][0] ),
    .A2(_03255_),
    .ZN(_03256_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07325_ (.A1(_03157_),
    .A2(_03255_),
    .B(_03256_),
    .ZN(_00551_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07326_ (.A1(\u_cpu.rf_ram.memory[49][1] ),
    .A2(_03255_),
    .ZN(_03257_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07327_ (.A1(_03161_),
    .A2(_03255_),
    .B(_03257_),
    .ZN(_00552_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07328_ (.A1(\u_cpu.rf_ram.memory[49][2] ),
    .A2(_03255_),
    .ZN(_03258_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07329_ (.A1(_03163_),
    .A2(_03255_),
    .B(_03258_),
    .ZN(_00553_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07330_ (.A1(\u_cpu.rf_ram.memory[49][3] ),
    .A2(_03255_),
    .ZN(_03259_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07331_ (.A1(_03165_),
    .A2(_03255_),
    .B(_03259_),
    .ZN(_00554_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07332_ (.A1(\u_cpu.rf_ram.memory[49][4] ),
    .A2(_03255_),
    .ZN(_03260_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07333_ (.A1(_03167_),
    .A2(_03255_),
    .B(_03260_),
    .ZN(_00555_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07334_ (.A1(\u_cpu.rf_ram.memory[49][5] ),
    .A2(_03255_),
    .ZN(_03261_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07335_ (.A1(_03169_),
    .A2(_03255_),
    .B(_03261_),
    .ZN(_00556_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07336_ (.A1(\u_cpu.rf_ram.memory[49][6] ),
    .A2(_03255_),
    .ZN(_03262_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07337_ (.A1(_03171_),
    .A2(_03255_),
    .B(_03262_),
    .ZN(_00557_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07338_ (.A1(\u_cpu.rf_ram.memory[49][7] ),
    .A2(_03255_),
    .ZN(_03263_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07339_ (.A1(_03173_),
    .A2(_03255_),
    .B(_03263_),
    .ZN(_00558_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07340_ (.A1(_02810_),
    .A2(_02832_),
    .ZN(_03264_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07341_ (.I(_03264_),
    .Z(_03265_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07342_ (.A1(\u_cpu.rf_ram.memory[136][0] ),
    .A2(_03265_),
    .ZN(_03266_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07343_ (.A1(_03157_),
    .A2(_03265_),
    .B(_03266_),
    .ZN(_00559_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07344_ (.A1(\u_cpu.rf_ram.memory[136][1] ),
    .A2(_03265_),
    .ZN(_03267_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07345_ (.A1(_03161_),
    .A2(_03265_),
    .B(_03267_),
    .ZN(_00560_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07346_ (.A1(\u_cpu.rf_ram.memory[136][2] ),
    .A2(_03265_),
    .ZN(_03268_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07347_ (.A1(_03163_),
    .A2(_03265_),
    .B(_03268_),
    .ZN(_00561_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07348_ (.A1(\u_cpu.rf_ram.memory[136][3] ),
    .A2(_03265_),
    .ZN(_03269_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07349_ (.A1(_03165_),
    .A2(_03265_),
    .B(_03269_),
    .ZN(_00562_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07350_ (.A1(\u_cpu.rf_ram.memory[136][4] ),
    .A2(_03265_),
    .ZN(_03270_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07351_ (.A1(_03167_),
    .A2(_03265_),
    .B(_03270_),
    .ZN(_00563_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07352_ (.A1(\u_cpu.rf_ram.memory[136][5] ),
    .A2(_03265_),
    .ZN(_03271_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07353_ (.A1(_03169_),
    .A2(_03265_),
    .B(_03271_),
    .ZN(_00564_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07354_ (.A1(\u_cpu.rf_ram.memory[136][6] ),
    .A2(_03265_),
    .ZN(_03272_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07355_ (.A1(_03171_),
    .A2(_03265_),
    .B(_03272_),
    .ZN(_00565_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07356_ (.A1(\u_cpu.rf_ram.memory[136][7] ),
    .A2(_03265_),
    .ZN(_03273_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07357_ (.A1(_03173_),
    .A2(_03265_),
    .B(_03273_),
    .ZN(_00566_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07358_ (.A1(_02602_),
    .A2(_02832_),
    .ZN(_03274_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07359_ (.I(_03274_),
    .Z(_03275_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07360_ (.A1(\u_cpu.rf_ram.memory[135][0] ),
    .A2(_03275_),
    .ZN(_03276_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07361_ (.A1(_03157_),
    .A2(_03275_),
    .B(_03276_),
    .ZN(_00567_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07362_ (.A1(\u_cpu.rf_ram.memory[135][1] ),
    .A2(_03275_),
    .ZN(_03277_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07363_ (.A1(_03161_),
    .A2(_03275_),
    .B(_03277_),
    .ZN(_00568_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07364_ (.A1(\u_cpu.rf_ram.memory[135][2] ),
    .A2(_03275_),
    .ZN(_03278_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07365_ (.A1(_03163_),
    .A2(_03275_),
    .B(_03278_),
    .ZN(_00569_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07366_ (.A1(\u_cpu.rf_ram.memory[135][3] ),
    .A2(_03275_),
    .ZN(_03279_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07367_ (.A1(_03165_),
    .A2(_03275_),
    .B(_03279_),
    .ZN(_00570_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07368_ (.A1(\u_cpu.rf_ram.memory[135][4] ),
    .A2(_03275_),
    .ZN(_03280_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07369_ (.A1(_03167_),
    .A2(_03275_),
    .B(_03280_),
    .ZN(_00571_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07370_ (.A1(\u_cpu.rf_ram.memory[135][5] ),
    .A2(_03275_),
    .ZN(_03281_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07371_ (.A1(_03169_),
    .A2(_03275_),
    .B(_03281_),
    .ZN(_00572_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07372_ (.A1(\u_cpu.rf_ram.memory[135][6] ),
    .A2(_03275_),
    .ZN(_03282_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07373_ (.A1(_03171_),
    .A2(_03275_),
    .B(_03282_),
    .ZN(_00573_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07374_ (.A1(\u_cpu.rf_ram.memory[135][7] ),
    .A2(_03275_),
    .ZN(_03283_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07375_ (.A1(_03173_),
    .A2(_03275_),
    .B(_03283_),
    .ZN(_00574_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07376_ (.A1(_02832_),
    .A2(_02893_),
    .ZN(_03284_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07377_ (.I(_03284_),
    .Z(_03285_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07378_ (.A1(\u_cpu.rf_ram.memory[134][0] ),
    .A2(_03285_),
    .ZN(_03286_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07379_ (.A1(_03157_),
    .A2(_03285_),
    .B(_03286_),
    .ZN(_00575_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07380_ (.A1(\u_cpu.rf_ram.memory[134][1] ),
    .A2(_03285_),
    .ZN(_03287_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07381_ (.A1(_03161_),
    .A2(_03285_),
    .B(_03287_),
    .ZN(_00576_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07382_ (.A1(\u_cpu.rf_ram.memory[134][2] ),
    .A2(_03285_),
    .ZN(_03288_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07383_ (.A1(_03163_),
    .A2(_03285_),
    .B(_03288_),
    .ZN(_00577_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07384_ (.A1(\u_cpu.rf_ram.memory[134][3] ),
    .A2(_03285_),
    .ZN(_03289_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07385_ (.A1(_03165_),
    .A2(_03285_),
    .B(_03289_),
    .ZN(_00578_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07386_ (.A1(\u_cpu.rf_ram.memory[134][4] ),
    .A2(_03285_),
    .ZN(_03290_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07387_ (.A1(_03167_),
    .A2(_03285_),
    .B(_03290_),
    .ZN(_00579_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07388_ (.A1(\u_cpu.rf_ram.memory[134][5] ),
    .A2(_03285_),
    .ZN(_03291_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07389_ (.A1(_03169_),
    .A2(_03285_),
    .B(_03291_),
    .ZN(_00580_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07390_ (.A1(\u_cpu.rf_ram.memory[134][6] ),
    .A2(_03285_),
    .ZN(_03292_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07391_ (.A1(_03171_),
    .A2(_03285_),
    .B(_03292_),
    .ZN(_00581_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07392_ (.A1(\u_cpu.rf_ram.memory[134][7] ),
    .A2(_03285_),
    .ZN(_03293_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07393_ (.A1(_03173_),
    .A2(_03285_),
    .B(_03293_),
    .ZN(_00582_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07394_ (.A1(_02524_),
    .A2(_02832_),
    .ZN(_03294_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07395_ (.I(_03294_),
    .Z(_03295_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07396_ (.A1(\u_cpu.rf_ram.memory[133][0] ),
    .A2(_03295_),
    .ZN(_03296_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07397_ (.A1(_03157_),
    .A2(_03295_),
    .B(_03296_),
    .ZN(_00583_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07398_ (.A1(\u_cpu.rf_ram.memory[133][1] ),
    .A2(_03295_),
    .ZN(_03297_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07399_ (.A1(_03161_),
    .A2(_03295_),
    .B(_03297_),
    .ZN(_00584_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07400_ (.A1(\u_cpu.rf_ram.memory[133][2] ),
    .A2(_03295_),
    .ZN(_03298_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07401_ (.A1(_03163_),
    .A2(_03295_),
    .B(_03298_),
    .ZN(_00585_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07402_ (.A1(\u_cpu.rf_ram.memory[133][3] ),
    .A2(_03295_),
    .ZN(_03299_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07403_ (.A1(_03165_),
    .A2(_03295_),
    .B(_03299_),
    .ZN(_00586_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07404_ (.A1(\u_cpu.rf_ram.memory[133][4] ),
    .A2(_03295_),
    .ZN(_03300_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07405_ (.A1(_03167_),
    .A2(_03295_),
    .B(_03300_),
    .ZN(_00587_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07406_ (.A1(\u_cpu.rf_ram.memory[133][5] ),
    .A2(_03295_),
    .ZN(_03301_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07407_ (.A1(_03169_),
    .A2(_03295_),
    .B(_03301_),
    .ZN(_00588_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07408_ (.A1(\u_cpu.rf_ram.memory[133][6] ),
    .A2(_03295_),
    .ZN(_03302_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07409_ (.A1(_03171_),
    .A2(_03295_),
    .B(_03302_),
    .ZN(_00589_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07410_ (.A1(\u_cpu.rf_ram.memory[133][7] ),
    .A2(_03295_),
    .ZN(_03303_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07411_ (.A1(_03173_),
    .A2(_03295_),
    .B(_03303_),
    .ZN(_00590_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07412_ (.A1(_02561_),
    .A2(_02832_),
    .ZN(_03304_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07413_ (.I(_03304_),
    .Z(_03305_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07414_ (.A1(\u_cpu.rf_ram.memory[132][0] ),
    .A2(_03305_),
    .ZN(_03306_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07415_ (.A1(_03157_),
    .A2(_03305_),
    .B(_03306_),
    .ZN(_00591_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07416_ (.A1(\u_cpu.rf_ram.memory[132][1] ),
    .A2(_03305_),
    .ZN(_03307_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07417_ (.A1(_03161_),
    .A2(_03305_),
    .B(_03307_),
    .ZN(_00592_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07418_ (.A1(\u_cpu.rf_ram.memory[132][2] ),
    .A2(_03305_),
    .ZN(_03308_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07419_ (.A1(_03163_),
    .A2(_03305_),
    .B(_03308_),
    .ZN(_00593_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07420_ (.A1(\u_cpu.rf_ram.memory[132][3] ),
    .A2(_03305_),
    .ZN(_03309_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07421_ (.A1(_03165_),
    .A2(_03305_),
    .B(_03309_),
    .ZN(_00594_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07422_ (.A1(\u_cpu.rf_ram.memory[132][4] ),
    .A2(_03305_),
    .ZN(_03310_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07423_ (.A1(_03167_),
    .A2(_03305_),
    .B(_03310_),
    .ZN(_00595_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07424_ (.A1(\u_cpu.rf_ram.memory[132][5] ),
    .A2(_03305_),
    .ZN(_03311_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07425_ (.A1(_03169_),
    .A2(_03305_),
    .B(_03311_),
    .ZN(_00596_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07426_ (.A1(\u_cpu.rf_ram.memory[132][6] ),
    .A2(_03305_),
    .ZN(_03312_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07427_ (.A1(_03171_),
    .A2(_03305_),
    .B(_03312_),
    .ZN(_00597_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07428_ (.A1(\u_cpu.rf_ram.memory[132][7] ),
    .A2(_03305_),
    .ZN(_03313_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07429_ (.A1(_03173_),
    .A2(_03305_),
    .B(_03313_),
    .ZN(_00598_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07430_ (.A1(_02682_),
    .A2(_02832_),
    .ZN(_03314_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07431_ (.I(_03314_),
    .Z(_03315_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07432_ (.A1(\u_cpu.rf_ram.memory[131][0] ),
    .A2(_03315_),
    .ZN(_03316_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07433_ (.A1(_03157_),
    .A2(_03315_),
    .B(_03316_),
    .ZN(_00599_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07434_ (.A1(\u_cpu.rf_ram.memory[131][1] ),
    .A2(_03315_),
    .ZN(_03317_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07435_ (.A1(_03161_),
    .A2(_03315_),
    .B(_03317_),
    .ZN(_00600_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07436_ (.A1(\u_cpu.rf_ram.memory[131][2] ),
    .A2(_03315_),
    .ZN(_03318_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07437_ (.A1(_03163_),
    .A2(_03315_),
    .B(_03318_),
    .ZN(_00601_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07438_ (.A1(\u_cpu.rf_ram.memory[131][3] ),
    .A2(_03315_),
    .ZN(_03319_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07439_ (.A1(_03165_),
    .A2(_03315_),
    .B(_03319_),
    .ZN(_00602_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07440_ (.A1(\u_cpu.rf_ram.memory[131][4] ),
    .A2(_03315_),
    .ZN(_03320_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07441_ (.A1(_03167_),
    .A2(_03315_),
    .B(_03320_),
    .ZN(_00603_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07442_ (.A1(\u_cpu.rf_ram.memory[131][5] ),
    .A2(_03315_),
    .ZN(_03321_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07443_ (.A1(_03169_),
    .A2(_03315_),
    .B(_03321_),
    .ZN(_00604_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07444_ (.A1(\u_cpu.rf_ram.memory[131][6] ),
    .A2(_03315_),
    .ZN(_03322_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07445_ (.A1(_03171_),
    .A2(_03315_),
    .B(_03322_),
    .ZN(_00605_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07446_ (.A1(\u_cpu.rf_ram.memory[131][7] ),
    .A2(_03315_),
    .ZN(_03323_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07447_ (.A1(_03173_),
    .A2(_03315_),
    .B(_03323_),
    .ZN(_00606_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07448_ (.A1(_02469_),
    .A2(_02832_),
    .ZN(_03324_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07449_ (.I(_03324_),
    .Z(_03325_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07450_ (.A1(\u_cpu.rf_ram.memory[130][0] ),
    .A2(_03325_),
    .ZN(_03326_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07451_ (.A1(_03157_),
    .A2(_03325_),
    .B(_03326_),
    .ZN(_00607_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07452_ (.A1(\u_cpu.rf_ram.memory[130][1] ),
    .A2(_03325_),
    .ZN(_03327_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07453_ (.A1(_03161_),
    .A2(_03325_),
    .B(_03327_),
    .ZN(_00608_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07454_ (.A1(\u_cpu.rf_ram.memory[130][2] ),
    .A2(_03325_),
    .ZN(_03328_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07455_ (.A1(_03163_),
    .A2(_03325_),
    .B(_03328_),
    .ZN(_00609_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07456_ (.A1(\u_cpu.rf_ram.memory[130][3] ),
    .A2(_03325_),
    .ZN(_03329_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07457_ (.A1(_03165_),
    .A2(_03325_),
    .B(_03329_),
    .ZN(_00610_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07458_ (.A1(\u_cpu.rf_ram.memory[130][4] ),
    .A2(_03325_),
    .ZN(_03330_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07459_ (.A1(_03167_),
    .A2(_03325_),
    .B(_03330_),
    .ZN(_00611_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07460_ (.A1(\u_cpu.rf_ram.memory[130][5] ),
    .A2(_03325_),
    .ZN(_03331_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07461_ (.A1(_03169_),
    .A2(_03325_),
    .B(_03331_),
    .ZN(_00612_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07462_ (.A1(\u_cpu.rf_ram.memory[130][6] ),
    .A2(_03325_),
    .ZN(_03332_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07463_ (.A1(_03171_),
    .A2(_03325_),
    .B(_03332_),
    .ZN(_00613_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07464_ (.A1(\u_cpu.rf_ram.memory[130][7] ),
    .A2(_03325_),
    .ZN(_03333_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07465_ (.A1(_03173_),
    .A2(_03325_),
    .B(_03333_),
    .ZN(_00614_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07466_ (.A1(_02577_),
    .A2(_02671_),
    .ZN(_03334_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07467_ (.I0(_02573_),
    .I1(\u_cpu.rf_ram.memory[12][0] ),
    .S(_03334_),
    .Z(_03335_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07468_ (.I(_03335_),
    .Z(_00615_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07469_ (.I0(_02581_),
    .I1(\u_cpu.rf_ram.memory[12][1] ),
    .S(_03334_),
    .Z(_03336_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07470_ (.I(_03336_),
    .Z(_00616_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07471_ (.I0(_02584_),
    .I1(\u_cpu.rf_ram.memory[12][2] ),
    .S(_03334_),
    .Z(_03337_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07472_ (.I(_03337_),
    .Z(_00617_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07473_ (.I0(_02587_),
    .I1(\u_cpu.rf_ram.memory[12][3] ),
    .S(_03334_),
    .Z(_03338_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07474_ (.I(_03338_),
    .Z(_00618_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07475_ (.I0(_02590_),
    .I1(\u_cpu.rf_ram.memory[12][4] ),
    .S(_03334_),
    .Z(_03339_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07476_ (.I(_03339_),
    .Z(_00619_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07477_ (.I0(_02593_),
    .I1(\u_cpu.rf_ram.memory[12][5] ),
    .S(_03334_),
    .Z(_03340_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07478_ (.I(_03340_),
    .Z(_00620_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07479_ (.I0(_02596_),
    .I1(\u_cpu.rf_ram.memory[12][6] ),
    .S(_03334_),
    .Z(_03341_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07480_ (.I(_03341_),
    .Z(_00621_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07481_ (.I0(_02599_),
    .I1(\u_cpu.rf_ram.memory[12][7] ),
    .S(_03334_),
    .Z(_03342_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07482_ (.I(_03342_),
    .Z(_00622_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07483_ (.I(_02481_),
    .Z(_03343_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07484_ (.A1(_02528_),
    .A2(_02893_),
    .ZN(_03344_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07485_ (.I(_03344_),
    .Z(_03345_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07486_ (.A1(\u_cpu.rf_ram.memory[22][0] ),
    .A2(_03345_),
    .ZN(_03346_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07487_ (.A1(_03343_),
    .A2(_03345_),
    .B(_03346_),
    .ZN(_00623_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07488_ (.I(_02486_),
    .Z(_03347_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07489_ (.A1(\u_cpu.rf_ram.memory[22][1] ),
    .A2(_03345_),
    .ZN(_03348_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07490_ (.A1(_03347_),
    .A2(_03345_),
    .B(_03348_),
    .ZN(_00624_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07491_ (.I(_02491_),
    .Z(_03349_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07492_ (.A1(\u_cpu.rf_ram.memory[22][2] ),
    .A2(_03345_),
    .ZN(_03350_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07493_ (.A1(_03349_),
    .A2(_03345_),
    .B(_03350_),
    .ZN(_00625_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07494_ (.I(_02496_),
    .Z(_03351_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07495_ (.A1(\u_cpu.rf_ram.memory[22][3] ),
    .A2(_03345_),
    .ZN(_03352_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07496_ (.A1(_03351_),
    .A2(_03345_),
    .B(_03352_),
    .ZN(_00626_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07497_ (.I(_02501_),
    .Z(_03353_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07498_ (.A1(\u_cpu.rf_ram.memory[22][4] ),
    .A2(_03345_),
    .ZN(_03354_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07499_ (.A1(_03353_),
    .A2(_03345_),
    .B(_03354_),
    .ZN(_00627_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07500_ (.I(_02506_),
    .Z(_03355_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07501_ (.A1(\u_cpu.rf_ram.memory[22][5] ),
    .A2(_03345_),
    .ZN(_03356_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07502_ (.A1(_03355_),
    .A2(_03345_),
    .B(_03356_),
    .ZN(_00628_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07503_ (.I(_02511_),
    .Z(_03357_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07504_ (.A1(\u_cpu.rf_ram.memory[22][6] ),
    .A2(_03345_),
    .ZN(_03358_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07505_ (.A1(_03357_),
    .A2(_03345_),
    .B(_03358_),
    .ZN(_00629_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07506_ (.I(_02516_),
    .Z(_03359_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07507_ (.A1(\u_cpu.rf_ram.memory[22][7] ),
    .A2(_03345_),
    .ZN(_03360_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07508_ (.A1(_03359_),
    .A2(_03345_),
    .B(_03360_),
    .ZN(_00630_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07509_ (.A1(_02612_),
    .A2(_02832_),
    .ZN(_03361_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07510_ (.I(_03361_),
    .Z(_03362_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07511_ (.A1(\u_cpu.rf_ram.memory[128][0] ),
    .A2(_03362_),
    .ZN(_03363_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07512_ (.A1(_03343_),
    .A2(_03362_),
    .B(_03363_),
    .ZN(_00631_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07513_ (.A1(\u_cpu.rf_ram.memory[128][1] ),
    .A2(_03362_),
    .ZN(_03364_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07514_ (.A1(_03347_),
    .A2(_03362_),
    .B(_03364_),
    .ZN(_00632_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07515_ (.A1(\u_cpu.rf_ram.memory[128][2] ),
    .A2(_03362_),
    .ZN(_03365_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07516_ (.A1(_03349_),
    .A2(_03362_),
    .B(_03365_),
    .ZN(_00633_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07517_ (.A1(\u_cpu.rf_ram.memory[128][3] ),
    .A2(_03362_),
    .ZN(_03366_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07518_ (.A1(_03351_),
    .A2(_03362_),
    .B(_03366_),
    .ZN(_00634_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07519_ (.A1(\u_cpu.rf_ram.memory[128][4] ),
    .A2(_03362_),
    .ZN(_03367_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07520_ (.A1(_03353_),
    .A2(_03362_),
    .B(_03367_),
    .ZN(_00635_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07521_ (.A1(\u_cpu.rf_ram.memory[128][5] ),
    .A2(_03362_),
    .ZN(_03368_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07522_ (.A1(_03355_),
    .A2(_03362_),
    .B(_03368_),
    .ZN(_00636_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07523_ (.A1(\u_cpu.rf_ram.memory[128][6] ),
    .A2(_03362_),
    .ZN(_03369_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07524_ (.A1(_03357_),
    .A2(_03362_),
    .B(_03369_),
    .ZN(_00637_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07525_ (.A1(\u_cpu.rf_ram.memory[128][7] ),
    .A2(_03362_),
    .ZN(_03370_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07526_ (.A1(_03359_),
    .A2(_03362_),
    .B(_03370_),
    .ZN(_00638_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07527_ (.A1(_02727_),
    .A2(_02821_),
    .ZN(_03371_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07528_ (.I(_03371_),
    .Z(_03372_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07529_ (.A1(\u_cpu.rf_ram.memory[127][0] ),
    .A2(_03372_),
    .ZN(_03373_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07530_ (.A1(_03343_),
    .A2(_03372_),
    .B(_03373_),
    .ZN(_00639_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07531_ (.A1(\u_cpu.rf_ram.memory[127][1] ),
    .A2(_03372_),
    .ZN(_03374_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07532_ (.A1(_03347_),
    .A2(_03372_),
    .B(_03374_),
    .ZN(_00640_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07533_ (.A1(\u_cpu.rf_ram.memory[127][2] ),
    .A2(_03372_),
    .ZN(_03375_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07534_ (.A1(_03349_),
    .A2(_03372_),
    .B(_03375_),
    .ZN(_00641_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07535_ (.A1(\u_cpu.rf_ram.memory[127][3] ),
    .A2(_03372_),
    .ZN(_03376_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07536_ (.A1(_03351_),
    .A2(_03372_),
    .B(_03376_),
    .ZN(_00642_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07537_ (.A1(\u_cpu.rf_ram.memory[127][4] ),
    .A2(_03372_),
    .ZN(_03377_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07538_ (.A1(_03353_),
    .A2(_03372_),
    .B(_03377_),
    .ZN(_00643_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07539_ (.A1(\u_cpu.rf_ram.memory[127][5] ),
    .A2(_03372_),
    .ZN(_03378_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07540_ (.A1(_03355_),
    .A2(_03372_),
    .B(_03378_),
    .ZN(_00644_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07541_ (.A1(\u_cpu.rf_ram.memory[127][6] ),
    .A2(_03372_),
    .ZN(_03379_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07542_ (.A1(_03357_),
    .A2(_03372_),
    .B(_03379_),
    .ZN(_00645_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07543_ (.A1(\u_cpu.rf_ram.memory[127][7] ),
    .A2(_03372_),
    .ZN(_03380_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07544_ (.A1(_03359_),
    .A2(_03372_),
    .B(_03380_),
    .ZN(_00646_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07545_ (.A1(_02625_),
    .A2(_02821_),
    .ZN(_03381_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07546_ (.I(_03381_),
    .Z(_03382_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07547_ (.A1(\u_cpu.rf_ram.memory[126][0] ),
    .A2(_03382_),
    .ZN(_03383_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07548_ (.A1(_03343_),
    .A2(_03382_),
    .B(_03383_),
    .ZN(_00647_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07549_ (.A1(\u_cpu.rf_ram.memory[126][1] ),
    .A2(_03382_),
    .ZN(_03384_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07550_ (.A1(_03347_),
    .A2(_03382_),
    .B(_03384_),
    .ZN(_00648_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07551_ (.A1(\u_cpu.rf_ram.memory[126][2] ),
    .A2(_03382_),
    .ZN(_03385_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07552_ (.A1(_03349_),
    .A2(_03382_),
    .B(_03385_),
    .ZN(_00649_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07553_ (.A1(\u_cpu.rf_ram.memory[126][3] ),
    .A2(_03382_),
    .ZN(_03386_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07554_ (.A1(_03351_),
    .A2(_03382_),
    .B(_03386_),
    .ZN(_00650_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07555_ (.A1(\u_cpu.rf_ram.memory[126][4] ),
    .A2(_03382_),
    .ZN(_03387_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07556_ (.A1(_03353_),
    .A2(_03382_),
    .B(_03387_),
    .ZN(_00651_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07557_ (.A1(\u_cpu.rf_ram.memory[126][5] ),
    .A2(_03382_),
    .ZN(_03388_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07558_ (.A1(_03355_),
    .A2(_03382_),
    .B(_03388_),
    .ZN(_00652_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07559_ (.A1(\u_cpu.rf_ram.memory[126][6] ),
    .A2(_03382_),
    .ZN(_03389_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07560_ (.A1(_03357_),
    .A2(_03382_),
    .B(_03389_),
    .ZN(_00653_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07561_ (.A1(\u_cpu.rf_ram.memory[126][7] ),
    .A2(_03382_),
    .ZN(_03390_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07562_ (.A1(_03359_),
    .A2(_03382_),
    .B(_03390_),
    .ZN(_00654_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07563_ (.A1(_02660_),
    .A2(_02821_),
    .ZN(_03391_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07564_ (.I(_03391_),
    .Z(_03392_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07565_ (.A1(\u_cpu.rf_ram.memory[125][0] ),
    .A2(_03392_),
    .ZN(_03393_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07566_ (.A1(_03343_),
    .A2(_03392_),
    .B(_03393_),
    .ZN(_00655_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07567_ (.A1(\u_cpu.rf_ram.memory[125][1] ),
    .A2(_03392_),
    .ZN(_03394_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07568_ (.A1(_03347_),
    .A2(_03392_),
    .B(_03394_),
    .ZN(_00656_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07569_ (.A1(\u_cpu.rf_ram.memory[125][2] ),
    .A2(_03392_),
    .ZN(_03395_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07570_ (.A1(_03349_),
    .A2(_03392_),
    .B(_03395_),
    .ZN(_00657_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07571_ (.A1(\u_cpu.rf_ram.memory[125][3] ),
    .A2(_03392_),
    .ZN(_03396_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07572_ (.A1(_03351_),
    .A2(_03392_),
    .B(_03396_),
    .ZN(_00658_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07573_ (.A1(\u_cpu.rf_ram.memory[125][4] ),
    .A2(_03392_),
    .ZN(_03397_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07574_ (.A1(_03353_),
    .A2(_03392_),
    .B(_03397_),
    .ZN(_00659_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07575_ (.A1(\u_cpu.rf_ram.memory[125][5] ),
    .A2(_03392_),
    .ZN(_03398_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07576_ (.A1(_03355_),
    .A2(_03392_),
    .B(_03398_),
    .ZN(_00660_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07577_ (.A1(\u_cpu.rf_ram.memory[125][6] ),
    .A2(_03392_),
    .ZN(_03399_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07578_ (.A1(_03357_),
    .A2(_03392_),
    .B(_03399_),
    .ZN(_00661_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07579_ (.A1(\u_cpu.rf_ram.memory[125][7] ),
    .A2(_03392_),
    .ZN(_03400_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07580_ (.A1(_03359_),
    .A2(_03392_),
    .B(_03400_),
    .ZN(_00662_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07581_ (.A1(_02671_),
    .A2(_02821_),
    .ZN(_03401_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07582_ (.I(_03401_),
    .Z(_03402_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07583_ (.A1(\u_cpu.rf_ram.memory[124][0] ),
    .A2(_03402_),
    .ZN(_03403_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07584_ (.A1(_03343_),
    .A2(_03402_),
    .B(_03403_),
    .ZN(_00663_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07585_ (.A1(\u_cpu.rf_ram.memory[124][1] ),
    .A2(_03402_),
    .ZN(_03404_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07586_ (.A1(_03347_),
    .A2(_03402_),
    .B(_03404_),
    .ZN(_00664_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07587_ (.A1(\u_cpu.rf_ram.memory[124][2] ),
    .A2(_03402_),
    .ZN(_03405_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07588_ (.A1(_03349_),
    .A2(_03402_),
    .B(_03405_),
    .ZN(_00665_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07589_ (.A1(\u_cpu.rf_ram.memory[124][3] ),
    .A2(_03402_),
    .ZN(_03406_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07590_ (.A1(_03351_),
    .A2(_03402_),
    .B(_03406_),
    .ZN(_00666_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07591_ (.A1(\u_cpu.rf_ram.memory[124][4] ),
    .A2(_03402_),
    .ZN(_03407_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07592_ (.A1(_03353_),
    .A2(_03402_),
    .B(_03407_),
    .ZN(_00667_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07593_ (.A1(\u_cpu.rf_ram.memory[124][5] ),
    .A2(_03402_),
    .ZN(_03408_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07594_ (.A1(_03355_),
    .A2(_03402_),
    .B(_03408_),
    .ZN(_00668_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07595_ (.A1(\u_cpu.rf_ram.memory[124][6] ),
    .A2(_03402_),
    .ZN(_03409_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07596_ (.A1(_03357_),
    .A2(_03402_),
    .B(_03409_),
    .ZN(_00669_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07597_ (.A1(\u_cpu.rf_ram.memory[124][7] ),
    .A2(_03402_),
    .ZN(_03410_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07598_ (.A1(_03359_),
    .A2(_03402_),
    .B(_03410_),
    .ZN(_00670_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07599_ (.A1(_02706_),
    .A2(_02821_),
    .ZN(_03411_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07600_ (.I(_03411_),
    .Z(_03412_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07601_ (.A1(\u_cpu.rf_ram.memory[123][0] ),
    .A2(_03412_),
    .ZN(_03413_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07602_ (.A1(_03343_),
    .A2(_03412_),
    .B(_03413_),
    .ZN(_00671_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07603_ (.A1(\u_cpu.rf_ram.memory[123][1] ),
    .A2(_03412_),
    .ZN(_03414_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07604_ (.A1(_03347_),
    .A2(_03412_),
    .B(_03414_),
    .ZN(_00672_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07605_ (.A1(\u_cpu.rf_ram.memory[123][2] ),
    .A2(_03412_),
    .ZN(_03415_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07606_ (.A1(_03349_),
    .A2(_03412_),
    .B(_03415_),
    .ZN(_00673_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07607_ (.A1(\u_cpu.rf_ram.memory[123][3] ),
    .A2(_03412_),
    .ZN(_03416_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07608_ (.A1(_03351_),
    .A2(_03412_),
    .B(_03416_),
    .ZN(_00674_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07609_ (.A1(\u_cpu.rf_ram.memory[123][4] ),
    .A2(_03412_),
    .ZN(_03417_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07610_ (.A1(_03353_),
    .A2(_03412_),
    .B(_03417_),
    .ZN(_00675_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07611_ (.A1(\u_cpu.rf_ram.memory[123][5] ),
    .A2(_03412_),
    .ZN(_03418_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07612_ (.A1(_03355_),
    .A2(_03412_),
    .B(_03418_),
    .ZN(_00676_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07613_ (.A1(\u_cpu.rf_ram.memory[123][6] ),
    .A2(_03412_),
    .ZN(_03419_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07614_ (.A1(_03357_),
    .A2(_03412_),
    .B(_03419_),
    .ZN(_00677_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07615_ (.A1(\u_cpu.rf_ram.memory[123][7] ),
    .A2(_03412_),
    .ZN(_03420_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07616_ (.A1(_03359_),
    .A2(_03412_),
    .B(_03420_),
    .ZN(_00678_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07617_ (.A1(_02639_),
    .A2(_02893_),
    .ZN(_03421_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07618_ (.I(_03421_),
    .Z(_03422_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07619_ (.A1(\u_cpu.rf_ram.memory[38][0] ),
    .A2(_03422_),
    .ZN(_03423_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07620_ (.A1(_03343_),
    .A2(_03422_),
    .B(_03423_),
    .ZN(_00679_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07621_ (.A1(\u_cpu.rf_ram.memory[38][1] ),
    .A2(_03422_),
    .ZN(_03424_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07622_ (.A1(_03347_),
    .A2(_03422_),
    .B(_03424_),
    .ZN(_00680_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07623_ (.A1(\u_cpu.rf_ram.memory[38][2] ),
    .A2(_03422_),
    .ZN(_03425_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07624_ (.A1(_03349_),
    .A2(_03422_),
    .B(_03425_),
    .ZN(_00681_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07625_ (.A1(\u_cpu.rf_ram.memory[38][3] ),
    .A2(_03422_),
    .ZN(_03426_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07626_ (.A1(_03351_),
    .A2(_03422_),
    .B(_03426_),
    .ZN(_00682_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07627_ (.A1(\u_cpu.rf_ram.memory[38][4] ),
    .A2(_03422_),
    .ZN(_03427_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07628_ (.A1(_03353_),
    .A2(_03422_),
    .B(_03427_),
    .ZN(_00683_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07629_ (.A1(\u_cpu.rf_ram.memory[38][5] ),
    .A2(_03422_),
    .ZN(_03428_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07630_ (.A1(_03355_),
    .A2(_03422_),
    .B(_03428_),
    .ZN(_00684_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07631_ (.A1(\u_cpu.rf_ram.memory[38][6] ),
    .A2(_03422_),
    .ZN(_03429_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07632_ (.A1(_03357_),
    .A2(_03422_),
    .B(_03429_),
    .ZN(_00685_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07633_ (.A1(\u_cpu.rf_ram.memory[38][7] ),
    .A2(_03422_),
    .ZN(_03430_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07634_ (.A1(_03359_),
    .A2(_03422_),
    .B(_03430_),
    .ZN(_00686_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07635_ (.A1(_02524_),
    .A2(_02639_),
    .ZN(_03431_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07636_ (.I(_03431_),
    .Z(_03432_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07637_ (.A1(\u_cpu.rf_ram.memory[37][0] ),
    .A2(_03432_),
    .ZN(_03433_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07638_ (.A1(_03343_),
    .A2(_03432_),
    .B(_03433_),
    .ZN(_00687_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07639_ (.A1(\u_cpu.rf_ram.memory[37][1] ),
    .A2(_03432_),
    .ZN(_03434_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07640_ (.A1(_03347_),
    .A2(_03432_),
    .B(_03434_),
    .ZN(_00688_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07641_ (.A1(\u_cpu.rf_ram.memory[37][2] ),
    .A2(_03432_),
    .ZN(_03435_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07642_ (.A1(_03349_),
    .A2(_03432_),
    .B(_03435_),
    .ZN(_00689_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07643_ (.A1(\u_cpu.rf_ram.memory[37][3] ),
    .A2(_03432_),
    .ZN(_03436_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07644_ (.A1(_03351_),
    .A2(_03432_),
    .B(_03436_),
    .ZN(_00690_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07645_ (.A1(\u_cpu.rf_ram.memory[37][4] ),
    .A2(_03432_),
    .ZN(_03437_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07646_ (.A1(_03353_),
    .A2(_03432_),
    .B(_03437_),
    .ZN(_00691_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07647_ (.A1(\u_cpu.rf_ram.memory[37][5] ),
    .A2(_03432_),
    .ZN(_03438_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07648_ (.A1(_03355_),
    .A2(_03432_),
    .B(_03438_),
    .ZN(_00692_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07649_ (.A1(\u_cpu.rf_ram.memory[37][6] ),
    .A2(_03432_),
    .ZN(_03439_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07650_ (.A1(_03357_),
    .A2(_03432_),
    .B(_03439_),
    .ZN(_00693_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07651_ (.A1(\u_cpu.rf_ram.memory[37][7] ),
    .A2(_03432_),
    .ZN(_03440_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07652_ (.A1(_03359_),
    .A2(_03432_),
    .B(_03440_),
    .ZN(_00694_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07653_ (.A1(_02561_),
    .A2(_02639_),
    .ZN(_03441_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07654_ (.I(_03441_),
    .Z(_03442_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07655_ (.A1(\u_cpu.rf_ram.memory[36][0] ),
    .A2(_03442_),
    .ZN(_03443_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07656_ (.A1(_03343_),
    .A2(_03442_),
    .B(_03443_),
    .ZN(_00695_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07657_ (.A1(\u_cpu.rf_ram.memory[36][1] ),
    .A2(_03442_),
    .ZN(_03444_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07658_ (.A1(_03347_),
    .A2(_03442_),
    .B(_03444_),
    .ZN(_00696_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07659_ (.A1(\u_cpu.rf_ram.memory[36][2] ),
    .A2(_03442_),
    .ZN(_03445_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07660_ (.A1(_03349_),
    .A2(_03442_),
    .B(_03445_),
    .ZN(_00697_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07661_ (.A1(\u_cpu.rf_ram.memory[36][3] ),
    .A2(_03442_),
    .ZN(_03446_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07662_ (.A1(_03351_),
    .A2(_03442_),
    .B(_03446_),
    .ZN(_00698_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07663_ (.A1(\u_cpu.rf_ram.memory[36][4] ),
    .A2(_03442_),
    .ZN(_03447_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07664_ (.A1(_03353_),
    .A2(_03442_),
    .B(_03447_),
    .ZN(_00699_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07665_ (.A1(\u_cpu.rf_ram.memory[36][5] ),
    .A2(_03442_),
    .ZN(_03448_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07666_ (.A1(_03355_),
    .A2(_03442_),
    .B(_03448_),
    .ZN(_00700_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07667_ (.A1(\u_cpu.rf_ram.memory[36][6] ),
    .A2(_03442_),
    .ZN(_03449_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07668_ (.A1(_03357_),
    .A2(_03442_),
    .B(_03449_),
    .ZN(_00701_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07669_ (.A1(\u_cpu.rf_ram.memory[36][7] ),
    .A2(_03442_),
    .ZN(_03450_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07670_ (.A1(_03359_),
    .A2(_03442_),
    .B(_03450_),
    .ZN(_00702_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07671_ (.A1(_02311_),
    .A2(_02773_),
    .ZN(_03451_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07672_ (.A1(_01428_),
    .A2(_03451_),
    .ZN(_03452_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07673_ (.I(_03452_),
    .Z(_00703_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07674_ (.A1(\u_cpu.cpu.state.o_cnt[2] ),
    .A2(\u_cpu.cpu.state.o_cnt_r[3] ),
    .ZN(_03453_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _07675_ (.A1(\u_cpu.cpu.state.o_cnt[2] ),
    .A2(\u_cpu.cpu.state.o_cnt_r[3] ),
    .Z(_03454_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _07676_ (.A1(_01428_),
    .A2(_03453_),
    .A3(_03454_),
    .ZN(_00704_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07677_ (.A1(\u_cpu.cpu.mem_bytecnt[0] ),
    .A2(_03454_),
    .B(_01429_),
    .ZN(_03455_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07678_ (.A1(\u_cpu.cpu.mem_bytecnt[0] ),
    .A2(_03454_),
    .B(_03455_),
    .ZN(_00705_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07679_ (.A1(\u_cpu.cpu.mem_bytecnt[0] ),
    .A2(_03454_),
    .ZN(_03456_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07680_ (.A1(\u_cpu.cpu.mem_bytecnt[1] ),
    .A2(_03456_),
    .Z(_03457_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07681_ (.A1(_01428_),
    .A2(_03457_),
    .ZN(_00706_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07682_ (.A1(_01428_),
    .A2(_02311_),
    .ZN(_03458_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07683_ (.A1(\u_cpu.cpu.state.o_cnt_r[3] ),
    .A2(_03458_),
    .ZN(_03459_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07684_ (.I(_02783_),
    .ZN(_03460_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07685_ (.A1(\u_cpu.rf_ram_if.rgnt ),
    .A2(_03460_),
    .B(_02433_),
    .C(_01429_),
    .ZN(_03461_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07686_ (.A1(_03459_),
    .A2(_03461_),
    .ZN(_00707_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _07687_ (.A1(_01429_),
    .A2(\u_cpu.cpu.state.o_cnt_r[0] ),
    .Z(_03462_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07688_ (.I(_03462_),
    .Z(_00708_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07689_ (.A1(_01428_),
    .A2(_02376_),
    .ZN(_00709_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _07690_ (.A1(_01429_),
    .A2(\u_cpu.cpu.state.o_cnt_r[2] ),
    .Z(_03463_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07691_ (.I(_03463_),
    .Z(_00710_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07692_ (.A1(_02475_),
    .A2(_02706_),
    .ZN(_03464_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07693_ (.I(_03464_),
    .Z(_03465_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07694_ (.A1(\u_cpu.rf_ram.memory[91][0] ),
    .A2(_03465_),
    .ZN(_03466_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07695_ (.A1(_03343_),
    .A2(_03465_),
    .B(_03466_),
    .ZN(_00711_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07696_ (.A1(\u_cpu.rf_ram.memory[91][1] ),
    .A2(_03465_),
    .ZN(_03467_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07697_ (.A1(_03347_),
    .A2(_03465_),
    .B(_03467_),
    .ZN(_00712_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07698_ (.A1(\u_cpu.rf_ram.memory[91][2] ),
    .A2(_03465_),
    .ZN(_03468_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07699_ (.A1(_03349_),
    .A2(_03465_),
    .B(_03468_),
    .ZN(_00713_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07700_ (.A1(\u_cpu.rf_ram.memory[91][3] ),
    .A2(_03465_),
    .ZN(_03469_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07701_ (.A1(_03351_),
    .A2(_03465_),
    .B(_03469_),
    .ZN(_00714_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07702_ (.A1(\u_cpu.rf_ram.memory[91][4] ),
    .A2(_03465_),
    .ZN(_03470_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07703_ (.A1(_03353_),
    .A2(_03465_),
    .B(_03470_),
    .ZN(_00715_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07704_ (.A1(\u_cpu.rf_ram.memory[91][5] ),
    .A2(_03465_),
    .ZN(_03471_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07705_ (.A1(_03355_),
    .A2(_03465_),
    .B(_03471_),
    .ZN(_00716_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07706_ (.A1(\u_cpu.rf_ram.memory[91][6] ),
    .A2(_03465_),
    .ZN(_03472_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07707_ (.A1(_03357_),
    .A2(_03465_),
    .B(_03472_),
    .ZN(_00717_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07708_ (.A1(\u_cpu.rf_ram.memory[91][7] ),
    .A2(_03465_),
    .ZN(_03473_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07709_ (.A1(_03359_),
    .A2(_03465_),
    .B(_03473_),
    .ZN(_00718_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07710_ (.A1(_02475_),
    .A2(_02638_),
    .ZN(_03474_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07711_ (.I(_03474_),
    .Z(_03475_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07712_ (.A1(\u_cpu.rf_ram.memory[90][0] ),
    .A2(_03475_),
    .ZN(_03476_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07713_ (.A1(_03343_),
    .A2(_03475_),
    .B(_03476_),
    .ZN(_00719_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07714_ (.A1(\u_cpu.rf_ram.memory[90][1] ),
    .A2(_03475_),
    .ZN(_03477_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07715_ (.A1(_03347_),
    .A2(_03475_),
    .B(_03477_),
    .ZN(_00720_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07716_ (.A1(\u_cpu.rf_ram.memory[90][2] ),
    .A2(_03475_),
    .ZN(_03478_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07717_ (.A1(_03349_),
    .A2(_03475_),
    .B(_03478_),
    .ZN(_00721_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07718_ (.A1(\u_cpu.rf_ram.memory[90][3] ),
    .A2(_03475_),
    .ZN(_03479_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07719_ (.A1(_03351_),
    .A2(_03475_),
    .B(_03479_),
    .ZN(_00722_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07720_ (.A1(\u_cpu.rf_ram.memory[90][4] ),
    .A2(_03475_),
    .ZN(_03480_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07721_ (.A1(_03353_),
    .A2(_03475_),
    .B(_03480_),
    .ZN(_00723_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07722_ (.A1(\u_cpu.rf_ram.memory[90][5] ),
    .A2(_03475_),
    .ZN(_03481_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07723_ (.A1(_03355_),
    .A2(_03475_),
    .B(_03481_),
    .ZN(_00724_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07724_ (.A1(\u_cpu.rf_ram.memory[90][6] ),
    .A2(_03475_),
    .ZN(_03482_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07725_ (.A1(_03357_),
    .A2(_03475_),
    .B(_03482_),
    .ZN(_00725_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07726_ (.A1(\u_cpu.rf_ram.memory[90][7] ),
    .A2(_03475_),
    .ZN(_03483_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07727_ (.A1(_03359_),
    .A2(_03475_),
    .B(_03483_),
    .ZN(_00726_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07728_ (.A1(_02432_),
    .A2(_02434_),
    .ZN(_03484_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07729_ (.A1(\u_cpu.cpu.state.genblk1.misalign_trap_sync_r ),
    .A2(_03458_),
    .ZN(_03485_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _07730_ (.A1(_01428_),
    .A2(_03451_),
    .A3(_03484_),
    .B(_03485_),
    .ZN(_00727_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07731_ (.A1(\u_cpu.cpu.ctrl.i_jump ),
    .A2(_03458_),
    .ZN(_03486_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07732_ (.A1(_02334_),
    .A2(_02364_),
    .ZN(_03487_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07733_ (.A1(_02309_),
    .A2(_03487_),
    .ZN(_03488_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _07734_ (.A1(_02325_),
    .A2(_03487_),
    .Z(_03489_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07735_ (.A1(_02328_),
    .A2(_03489_),
    .Z(_03490_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _07736_ (.A1(_03488_),
    .A2(_03490_),
    .Z(_03491_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07737_ (.A1(_01408_),
    .A2(_02332_),
    .B1(_03488_),
    .B2(_03490_),
    .ZN(_03492_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _07738_ (.A1(_02355_),
    .A2(_02356_),
    .B(_01369_),
    .C(_01370_),
    .ZN(_03493_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07739_ (.A1(_03491_),
    .A2(_03492_),
    .B1(_03493_),
    .B2(_02359_),
    .ZN(_03494_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07740_ (.A1(_02333_),
    .A2(_03494_),
    .Z(_03495_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07741_ (.A1(_02313_),
    .A2(_03495_),
    .B(_00703_),
    .C(_01374_),
    .ZN(_03496_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07742_ (.A1(_03486_),
    .A2(_03496_),
    .ZN(_00729_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _07743_ (.A1(\u_cpu.cpu.mem_bytecnt[1] ),
    .A2(_02395_),
    .A3(_00710_),
    .Z(_03497_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07744_ (.I(_03497_),
    .Z(_00730_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07745_ (.A1(\u_cpu.cpu.state.init_done ),
    .A2(_03458_),
    .ZN(_03498_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07746_ (.A1(_01428_),
    .A2(_03451_),
    .B(_03498_),
    .ZN(_00731_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07747_ (.A1(_02475_),
    .A2(_02671_),
    .ZN(_03499_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07748_ (.I(_03499_),
    .Z(_03500_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07749_ (.A1(\u_cpu.rf_ram.memory[92][0] ),
    .A2(_03500_),
    .ZN(_03501_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07750_ (.A1(_03343_),
    .A2(_03500_),
    .B(_03501_),
    .ZN(_00732_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07751_ (.A1(\u_cpu.rf_ram.memory[92][1] ),
    .A2(_03500_),
    .ZN(_03502_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07752_ (.A1(_03347_),
    .A2(_03500_),
    .B(_03502_),
    .ZN(_00733_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07753_ (.A1(\u_cpu.rf_ram.memory[92][2] ),
    .A2(_03500_),
    .ZN(_03503_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07754_ (.A1(_03349_),
    .A2(_03500_),
    .B(_03503_),
    .ZN(_00734_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07755_ (.A1(\u_cpu.rf_ram.memory[92][3] ),
    .A2(_03500_),
    .ZN(_03504_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07756_ (.A1(_03351_),
    .A2(_03500_),
    .B(_03504_),
    .ZN(_00735_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07757_ (.A1(\u_cpu.rf_ram.memory[92][4] ),
    .A2(_03500_),
    .ZN(_03505_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07758_ (.A1(_03353_),
    .A2(_03500_),
    .B(_03505_),
    .ZN(_00736_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07759_ (.A1(\u_cpu.rf_ram.memory[92][5] ),
    .A2(_03500_),
    .ZN(_03506_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07760_ (.A1(_03355_),
    .A2(_03500_),
    .B(_03506_),
    .ZN(_00737_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07761_ (.A1(\u_cpu.rf_ram.memory[92][6] ),
    .A2(_03500_),
    .ZN(_03507_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07762_ (.A1(_03357_),
    .A2(_03500_),
    .B(_03507_),
    .ZN(_00738_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07763_ (.A1(\u_cpu.rf_ram.memory[92][7] ),
    .A2(_03500_),
    .ZN(_03508_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07764_ (.A1(_03359_),
    .A2(_03500_),
    .B(_03508_),
    .ZN(_00739_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07765_ (.A1(_02639_),
    .A2(_02682_),
    .ZN(_03509_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07766_ (.I(_03509_),
    .Z(_03510_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07767_ (.A1(\u_cpu.rf_ram.memory[35][0] ),
    .A2(_03510_),
    .ZN(_03511_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07768_ (.A1(_03343_),
    .A2(_03510_),
    .B(_03511_),
    .ZN(_00740_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07769_ (.A1(\u_cpu.rf_ram.memory[35][1] ),
    .A2(_03510_),
    .ZN(_03512_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07770_ (.A1(_03347_),
    .A2(_03510_),
    .B(_03512_),
    .ZN(_00741_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07771_ (.A1(\u_cpu.rf_ram.memory[35][2] ),
    .A2(_03510_),
    .ZN(_03513_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07772_ (.A1(_03349_),
    .A2(_03510_),
    .B(_03513_),
    .ZN(_00742_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07773_ (.A1(\u_cpu.rf_ram.memory[35][3] ),
    .A2(_03510_),
    .ZN(_03514_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07774_ (.A1(_03351_),
    .A2(_03510_),
    .B(_03514_),
    .ZN(_00743_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07775_ (.A1(\u_cpu.rf_ram.memory[35][4] ),
    .A2(_03510_),
    .ZN(_03515_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07776_ (.A1(_03353_),
    .A2(_03510_),
    .B(_03515_),
    .ZN(_00744_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07777_ (.A1(\u_cpu.rf_ram.memory[35][5] ),
    .A2(_03510_),
    .ZN(_03516_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07778_ (.A1(_03355_),
    .A2(_03510_),
    .B(_03516_),
    .ZN(_00745_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07779_ (.A1(\u_cpu.rf_ram.memory[35][6] ),
    .A2(_03510_),
    .ZN(_03517_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07780_ (.A1(_03357_),
    .A2(_03510_),
    .B(_03517_),
    .ZN(_00746_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07781_ (.A1(\u_cpu.rf_ram.memory[35][7] ),
    .A2(_03510_),
    .ZN(_03518_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07782_ (.A1(_03359_),
    .A2(_03510_),
    .B(_03518_),
    .ZN(_00747_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07783_ (.A1(_02469_),
    .A2(_02639_),
    .ZN(_03519_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07784_ (.I(_03519_),
    .Z(_03520_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07785_ (.A1(\u_cpu.rf_ram.memory[34][0] ),
    .A2(_03520_),
    .ZN(_03521_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07786_ (.A1(_03343_),
    .A2(_03520_),
    .B(_03521_),
    .ZN(_00748_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07787_ (.A1(\u_cpu.rf_ram.memory[34][1] ),
    .A2(_03520_),
    .ZN(_03522_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07788_ (.A1(_03347_),
    .A2(_03520_),
    .B(_03522_),
    .ZN(_00749_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07789_ (.A1(\u_cpu.rf_ram.memory[34][2] ),
    .A2(_03520_),
    .ZN(_03523_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07790_ (.A1(_03349_),
    .A2(_03520_),
    .B(_03523_),
    .ZN(_00750_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07791_ (.A1(\u_cpu.rf_ram.memory[34][3] ),
    .A2(_03520_),
    .ZN(_03524_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07792_ (.A1(_03351_),
    .A2(_03520_),
    .B(_03524_),
    .ZN(_00751_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07793_ (.A1(\u_cpu.rf_ram.memory[34][4] ),
    .A2(_03520_),
    .ZN(_03525_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07794_ (.A1(_03353_),
    .A2(_03520_),
    .B(_03525_),
    .ZN(_00752_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07795_ (.A1(\u_cpu.rf_ram.memory[34][5] ),
    .A2(_03520_),
    .ZN(_03526_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07796_ (.A1(_03355_),
    .A2(_03520_),
    .B(_03526_),
    .ZN(_00753_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07797_ (.A1(\u_cpu.rf_ram.memory[34][6] ),
    .A2(_03520_),
    .ZN(_03527_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07798_ (.A1(_03357_),
    .A2(_03520_),
    .B(_03527_),
    .ZN(_00754_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07799_ (.A1(\u_cpu.rf_ram.memory[34][7] ),
    .A2(_03520_),
    .ZN(_03528_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07800_ (.A1(_03359_),
    .A2(_03520_),
    .B(_03528_),
    .ZN(_00755_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07801_ (.A1(_02524_),
    .A2(_02821_),
    .ZN(_03529_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07802_ (.I(_03529_),
    .Z(_03530_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07803_ (.A1(\u_cpu.rf_ram.memory[117][0] ),
    .A2(_03530_),
    .ZN(_03531_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07804_ (.A1(_03343_),
    .A2(_03530_),
    .B(_03531_),
    .ZN(_00756_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07805_ (.A1(\u_cpu.rf_ram.memory[117][1] ),
    .A2(_03530_),
    .ZN(_03532_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07806_ (.A1(_03347_),
    .A2(_03530_),
    .B(_03532_),
    .ZN(_00757_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07807_ (.A1(\u_cpu.rf_ram.memory[117][2] ),
    .A2(_03530_),
    .ZN(_03533_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07808_ (.A1(_03349_),
    .A2(_03530_),
    .B(_03533_),
    .ZN(_00758_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07809_ (.A1(\u_cpu.rf_ram.memory[117][3] ),
    .A2(_03530_),
    .ZN(_03534_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07810_ (.A1(_03351_),
    .A2(_03530_),
    .B(_03534_),
    .ZN(_00759_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07811_ (.A1(\u_cpu.rf_ram.memory[117][4] ),
    .A2(_03530_),
    .ZN(_03535_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07812_ (.A1(_03353_),
    .A2(_03530_),
    .B(_03535_),
    .ZN(_00760_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07813_ (.A1(\u_cpu.rf_ram.memory[117][5] ),
    .A2(_03530_),
    .ZN(_03536_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07814_ (.A1(_03355_),
    .A2(_03530_),
    .B(_03536_),
    .ZN(_00761_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07815_ (.A1(\u_cpu.rf_ram.memory[117][6] ),
    .A2(_03530_),
    .ZN(_03537_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07816_ (.A1(_03357_),
    .A2(_03530_),
    .B(_03537_),
    .ZN(_00762_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07817_ (.A1(\u_cpu.rf_ram.memory[117][7] ),
    .A2(_03530_),
    .ZN(_03538_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07818_ (.A1(_03359_),
    .A2(_03530_),
    .B(_03538_),
    .ZN(_00763_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07819_ (.I(_02481_),
    .Z(_03539_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07820_ (.A1(_02810_),
    .A2(_02821_),
    .ZN(_03540_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07821_ (.I(_03540_),
    .Z(_03541_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07822_ (.A1(\u_cpu.rf_ram.memory[120][0] ),
    .A2(_03541_),
    .ZN(_03542_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07823_ (.A1(_03539_),
    .A2(_03541_),
    .B(_03542_),
    .ZN(_00764_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07824_ (.I(_02486_),
    .Z(_03543_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07825_ (.A1(\u_cpu.rf_ram.memory[120][1] ),
    .A2(_03541_),
    .ZN(_03544_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07826_ (.A1(_03543_),
    .A2(_03541_),
    .B(_03544_),
    .ZN(_00765_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07827_ (.I(_02491_),
    .Z(_03545_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07828_ (.A1(\u_cpu.rf_ram.memory[120][2] ),
    .A2(_03541_),
    .ZN(_03546_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07829_ (.A1(_03545_),
    .A2(_03541_),
    .B(_03546_),
    .ZN(_00766_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07830_ (.I(_02496_),
    .Z(_03547_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07831_ (.A1(\u_cpu.rf_ram.memory[120][3] ),
    .A2(_03541_),
    .ZN(_03548_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07832_ (.A1(_03547_),
    .A2(_03541_),
    .B(_03548_),
    .ZN(_00767_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07833_ (.I(_02501_),
    .Z(_03549_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07834_ (.A1(\u_cpu.rf_ram.memory[120][4] ),
    .A2(_03541_),
    .ZN(_03550_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07835_ (.A1(_03549_),
    .A2(_03541_),
    .B(_03550_),
    .ZN(_00768_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07836_ (.I(_02506_),
    .Z(_03551_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07837_ (.A1(\u_cpu.rf_ram.memory[120][5] ),
    .A2(_03541_),
    .ZN(_03552_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07838_ (.A1(_03551_),
    .A2(_03541_),
    .B(_03552_),
    .ZN(_00769_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07839_ (.I(_02511_),
    .Z(_03553_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07840_ (.A1(\u_cpu.rf_ram.memory[120][6] ),
    .A2(_03541_),
    .ZN(_03554_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07841_ (.A1(_03553_),
    .A2(_03541_),
    .B(_03554_),
    .ZN(_00770_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07842_ (.I(_02516_),
    .Z(_03555_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07843_ (.A1(\u_cpu.rf_ram.memory[120][7] ),
    .A2(_03541_),
    .ZN(_03556_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07844_ (.A1(_03555_),
    .A2(_03541_),
    .B(_03556_),
    .ZN(_00771_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07845_ (.A1(_02821_),
    .A2(_02893_),
    .ZN(_03557_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07846_ (.I(_03557_),
    .Z(_03558_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07847_ (.A1(\u_cpu.rf_ram.memory[118][0] ),
    .A2(_03558_),
    .ZN(_03559_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07848_ (.A1(_03539_),
    .A2(_03558_),
    .B(_03559_),
    .ZN(_00772_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07849_ (.A1(\u_cpu.rf_ram.memory[118][1] ),
    .A2(_03558_),
    .ZN(_03560_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07850_ (.A1(_03543_),
    .A2(_03558_),
    .B(_03560_),
    .ZN(_00773_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07851_ (.A1(\u_cpu.rf_ram.memory[118][2] ),
    .A2(_03558_),
    .ZN(_03561_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07852_ (.A1(_03545_),
    .A2(_03558_),
    .B(_03561_),
    .ZN(_00774_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07853_ (.A1(\u_cpu.rf_ram.memory[118][3] ),
    .A2(_03558_),
    .ZN(_03562_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07854_ (.A1(_03547_),
    .A2(_03558_),
    .B(_03562_),
    .ZN(_00775_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07855_ (.A1(\u_cpu.rf_ram.memory[118][4] ),
    .A2(_03558_),
    .ZN(_03563_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07856_ (.A1(_03549_),
    .A2(_03558_),
    .B(_03563_),
    .ZN(_00776_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07857_ (.A1(\u_cpu.rf_ram.memory[118][5] ),
    .A2(_03558_),
    .ZN(_03564_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07858_ (.A1(_03551_),
    .A2(_03558_),
    .B(_03564_),
    .ZN(_00777_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07859_ (.A1(\u_cpu.rf_ram.memory[118][6] ),
    .A2(_03558_),
    .ZN(_03565_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07860_ (.A1(_03553_),
    .A2(_03558_),
    .B(_03565_),
    .ZN(_00778_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07861_ (.A1(\u_cpu.rf_ram.memory[118][7] ),
    .A2(_03558_),
    .ZN(_03566_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07862_ (.A1(_03555_),
    .A2(_03558_),
    .B(_03566_),
    .ZN(_00779_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07863_ (.A1(_02695_),
    .A2(_02821_),
    .ZN(_03567_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07864_ (.I(_03567_),
    .Z(_03568_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07865_ (.A1(\u_cpu.rf_ram.memory[121][0] ),
    .A2(_03568_),
    .ZN(_03569_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07866_ (.A1(_03539_),
    .A2(_03568_),
    .B(_03569_),
    .ZN(_00780_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07867_ (.A1(\u_cpu.rf_ram.memory[121][1] ),
    .A2(_03568_),
    .ZN(_03570_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07868_ (.A1(_03543_),
    .A2(_03568_),
    .B(_03570_),
    .ZN(_00781_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07869_ (.A1(\u_cpu.rf_ram.memory[121][2] ),
    .A2(_03568_),
    .ZN(_03571_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07870_ (.A1(_03545_),
    .A2(_03568_),
    .B(_03571_),
    .ZN(_00782_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07871_ (.A1(\u_cpu.rf_ram.memory[121][3] ),
    .A2(_03568_),
    .ZN(_03572_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07872_ (.A1(_03547_),
    .A2(_03568_),
    .B(_03572_),
    .ZN(_00783_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07873_ (.A1(\u_cpu.rf_ram.memory[121][4] ),
    .A2(_03568_),
    .ZN(_03573_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07874_ (.A1(_03549_),
    .A2(_03568_),
    .B(_03573_),
    .ZN(_00784_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07875_ (.A1(\u_cpu.rf_ram.memory[121][5] ),
    .A2(_03568_),
    .ZN(_03574_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07876_ (.A1(_03551_),
    .A2(_03568_),
    .B(_03574_),
    .ZN(_00785_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07877_ (.A1(\u_cpu.rf_ram.memory[121][6] ),
    .A2(_03568_),
    .ZN(_03575_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07878_ (.A1(_03553_),
    .A2(_03568_),
    .B(_03575_),
    .ZN(_00786_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07879_ (.A1(\u_cpu.rf_ram.memory[121][7] ),
    .A2(_03568_),
    .ZN(_03576_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07880_ (.A1(_03555_),
    .A2(_03568_),
    .B(_03576_),
    .ZN(_00787_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07881_ (.A1(_02577_),
    .A2(_02810_),
    .ZN(_03577_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07882_ (.I0(_02573_),
    .I1(\u_cpu.rf_ram.memory[8][0] ),
    .S(_03577_),
    .Z(_03578_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07883_ (.I(_03578_),
    .Z(_00788_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07884_ (.I0(_02581_),
    .I1(\u_cpu.rf_ram.memory[8][1] ),
    .S(_03577_),
    .Z(_03579_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07885_ (.I(_03579_),
    .Z(_00789_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07886_ (.I0(_02584_),
    .I1(\u_cpu.rf_ram.memory[8][2] ),
    .S(_03577_),
    .Z(_03580_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07887_ (.I(_03580_),
    .Z(_00790_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07888_ (.I0(_02587_),
    .I1(\u_cpu.rf_ram.memory[8][3] ),
    .S(_03577_),
    .Z(_03581_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07889_ (.I(_03581_),
    .Z(_00791_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07890_ (.I0(_02590_),
    .I1(\u_cpu.rf_ram.memory[8][4] ),
    .S(_03577_),
    .Z(_03582_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07891_ (.I(_03582_),
    .Z(_00792_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07892_ (.I0(_02593_),
    .I1(\u_cpu.rf_ram.memory[8][5] ),
    .S(_03577_),
    .Z(_03583_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07893_ (.I(_03583_),
    .Z(_00793_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07894_ (.I0(_02596_),
    .I1(\u_cpu.rf_ram.memory[8][6] ),
    .S(_03577_),
    .Z(_03584_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07895_ (.I(_03584_),
    .Z(_00794_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07896_ (.I0(_02599_),
    .I1(\u_cpu.rf_ram.memory[8][7] ),
    .S(_03577_),
    .Z(_03585_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07897_ (.I(_03585_),
    .Z(_00795_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07898_ (.A1(_02577_),
    .A2(_02706_),
    .ZN(_03586_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07899_ (.I0(_02573_),
    .I1(\u_cpu.rf_ram.memory[11][0] ),
    .S(_03586_),
    .Z(_03587_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07900_ (.I(_03587_),
    .Z(_00796_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07901_ (.I0(_02581_),
    .I1(\u_cpu.rf_ram.memory[11][1] ),
    .S(_03586_),
    .Z(_03588_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07902_ (.I(_03588_),
    .Z(_00797_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07903_ (.I0(_02584_),
    .I1(\u_cpu.rf_ram.memory[11][2] ),
    .S(_03586_),
    .Z(_03589_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07904_ (.I(_03589_),
    .Z(_00798_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07905_ (.I0(_02587_),
    .I1(\u_cpu.rf_ram.memory[11][3] ),
    .S(_03586_),
    .Z(_03590_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07906_ (.I(_03590_),
    .Z(_00799_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07907_ (.I0(_02590_),
    .I1(\u_cpu.rf_ram.memory[11][4] ),
    .S(_03586_),
    .Z(_03591_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07908_ (.I(_03591_),
    .Z(_00800_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07909_ (.I0(_02593_),
    .I1(\u_cpu.rf_ram.memory[11][5] ),
    .S(_03586_),
    .Z(_03592_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07910_ (.I(_03592_),
    .Z(_00801_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07911_ (.I0(_02596_),
    .I1(\u_cpu.rf_ram.memory[11][6] ),
    .S(_03586_),
    .Z(_03593_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07912_ (.I(_03593_),
    .Z(_00802_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07913_ (.I0(_02599_),
    .I1(\u_cpu.rf_ram.memory[11][7] ),
    .S(_03586_),
    .Z(_03594_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07914_ (.I(_03594_),
    .Z(_00803_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07915_ (.A1(_02612_),
    .A2(_02821_),
    .ZN(_03595_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07916_ (.I(_03595_),
    .Z(_03596_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07917_ (.A1(\u_cpu.rf_ram.memory[112][0] ),
    .A2(_03596_),
    .ZN(_03597_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07918_ (.A1(_03539_),
    .A2(_03596_),
    .B(_03597_),
    .ZN(_00804_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07919_ (.A1(\u_cpu.rf_ram.memory[112][1] ),
    .A2(_03596_),
    .ZN(_03598_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07920_ (.A1(_03543_),
    .A2(_03596_),
    .B(_03598_),
    .ZN(_00805_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07921_ (.A1(\u_cpu.rf_ram.memory[112][2] ),
    .A2(_03596_),
    .ZN(_03599_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07922_ (.A1(_03545_),
    .A2(_03596_),
    .B(_03599_),
    .ZN(_00806_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07923_ (.A1(\u_cpu.rf_ram.memory[112][3] ),
    .A2(_03596_),
    .ZN(_03600_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07924_ (.A1(_03547_),
    .A2(_03596_),
    .B(_03600_),
    .ZN(_00807_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07925_ (.A1(\u_cpu.rf_ram.memory[112][4] ),
    .A2(_03596_),
    .ZN(_03601_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07926_ (.A1(_03549_),
    .A2(_03596_),
    .B(_03601_),
    .ZN(_00808_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07927_ (.A1(\u_cpu.rf_ram.memory[112][5] ),
    .A2(_03596_),
    .ZN(_03602_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07928_ (.A1(_03551_),
    .A2(_03596_),
    .B(_03602_),
    .ZN(_00809_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07929_ (.A1(\u_cpu.rf_ram.memory[112][6] ),
    .A2(_03596_),
    .ZN(_03603_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07930_ (.A1(_03553_),
    .A2(_03596_),
    .B(_03603_),
    .ZN(_00810_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07931_ (.A1(\u_cpu.rf_ram.memory[112][7] ),
    .A2(_03596_),
    .ZN(_03604_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07932_ (.A1(_03555_),
    .A2(_03596_),
    .B(_03604_),
    .ZN(_00811_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07933_ (.A1(_02638_),
    .A2(_02821_),
    .ZN(_03605_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07934_ (.I(_03605_),
    .Z(_03606_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07935_ (.A1(\u_cpu.rf_ram.memory[122][0] ),
    .A2(_03606_),
    .ZN(_03607_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07936_ (.A1(_03539_),
    .A2(_03606_),
    .B(_03607_),
    .ZN(_00812_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07937_ (.A1(\u_cpu.rf_ram.memory[122][1] ),
    .A2(_03606_),
    .ZN(_03608_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07938_ (.A1(_03543_),
    .A2(_03606_),
    .B(_03608_),
    .ZN(_00813_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07939_ (.A1(\u_cpu.rf_ram.memory[122][2] ),
    .A2(_03606_),
    .ZN(_03609_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07940_ (.A1(_03545_),
    .A2(_03606_),
    .B(_03609_),
    .ZN(_00814_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07941_ (.A1(\u_cpu.rf_ram.memory[122][3] ),
    .A2(_03606_),
    .ZN(_03610_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07942_ (.A1(_03547_),
    .A2(_03606_),
    .B(_03610_),
    .ZN(_00815_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07943_ (.A1(\u_cpu.rf_ram.memory[122][4] ),
    .A2(_03606_),
    .ZN(_03611_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07944_ (.A1(_03549_),
    .A2(_03606_),
    .B(_03611_),
    .ZN(_00816_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07945_ (.A1(\u_cpu.rf_ram.memory[122][5] ),
    .A2(_03606_),
    .ZN(_03612_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07946_ (.A1(_03551_),
    .A2(_03606_),
    .B(_03612_),
    .ZN(_00817_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07947_ (.A1(\u_cpu.rf_ram.memory[122][6] ),
    .A2(_03606_),
    .ZN(_03613_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07948_ (.A1(_03553_),
    .A2(_03606_),
    .B(_03613_),
    .ZN(_00818_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07949_ (.A1(\u_cpu.rf_ram.memory[122][7] ),
    .A2(_03606_),
    .ZN(_03614_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07950_ (.A1(_03555_),
    .A2(_03606_),
    .B(_03614_),
    .ZN(_00819_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07951_ (.A1(_02682_),
    .A2(_02821_),
    .ZN(_03615_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07952_ (.I(_03615_),
    .Z(_03616_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07953_ (.A1(\u_cpu.rf_ram.memory[115][0] ),
    .A2(_03616_),
    .ZN(_03617_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07954_ (.A1(_03539_),
    .A2(_03616_),
    .B(_03617_),
    .ZN(_00820_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07955_ (.A1(\u_cpu.rf_ram.memory[115][1] ),
    .A2(_03616_),
    .ZN(_03618_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07956_ (.A1(_03543_),
    .A2(_03616_),
    .B(_03618_),
    .ZN(_00821_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07957_ (.A1(\u_cpu.rf_ram.memory[115][2] ),
    .A2(_03616_),
    .ZN(_03619_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07958_ (.A1(_03545_),
    .A2(_03616_),
    .B(_03619_),
    .ZN(_00822_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07959_ (.A1(\u_cpu.rf_ram.memory[115][3] ),
    .A2(_03616_),
    .ZN(_03620_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07960_ (.A1(_03547_),
    .A2(_03616_),
    .B(_03620_),
    .ZN(_00823_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07961_ (.A1(\u_cpu.rf_ram.memory[115][4] ),
    .A2(_03616_),
    .ZN(_03621_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07962_ (.A1(_03549_),
    .A2(_03616_),
    .B(_03621_),
    .ZN(_00824_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07963_ (.A1(\u_cpu.rf_ram.memory[115][5] ),
    .A2(_03616_),
    .ZN(_03622_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07964_ (.A1(_03551_),
    .A2(_03616_),
    .B(_03622_),
    .ZN(_00825_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07965_ (.A1(\u_cpu.rf_ram.memory[115][6] ),
    .A2(_03616_),
    .ZN(_03623_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07966_ (.A1(_03553_),
    .A2(_03616_),
    .B(_03623_),
    .ZN(_00826_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07967_ (.A1(\u_cpu.rf_ram.memory[115][7] ),
    .A2(_03616_),
    .ZN(_03624_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07968_ (.A1(_03555_),
    .A2(_03616_),
    .B(_03624_),
    .ZN(_00827_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07969_ (.A1(_02561_),
    .A2(_02821_),
    .ZN(_03625_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07970_ (.I(_03625_),
    .Z(_03626_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07971_ (.A1(\u_cpu.rf_ram.memory[116][0] ),
    .A2(_03626_),
    .ZN(_03627_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07972_ (.A1(_03539_),
    .A2(_03626_),
    .B(_03627_),
    .ZN(_00828_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07973_ (.A1(\u_cpu.rf_ram.memory[116][1] ),
    .A2(_03626_),
    .ZN(_03628_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07974_ (.A1(_03543_),
    .A2(_03626_),
    .B(_03628_),
    .ZN(_00829_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07975_ (.A1(\u_cpu.rf_ram.memory[116][2] ),
    .A2(_03626_),
    .ZN(_03629_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07976_ (.A1(_03545_),
    .A2(_03626_),
    .B(_03629_),
    .ZN(_00830_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07977_ (.A1(\u_cpu.rf_ram.memory[116][3] ),
    .A2(_03626_),
    .ZN(_03630_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07978_ (.A1(_03547_),
    .A2(_03626_),
    .B(_03630_),
    .ZN(_00831_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07979_ (.A1(\u_cpu.rf_ram.memory[116][4] ),
    .A2(_03626_),
    .ZN(_03631_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07980_ (.A1(_03549_),
    .A2(_03626_),
    .B(_03631_),
    .ZN(_00832_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07981_ (.A1(\u_cpu.rf_ram.memory[116][5] ),
    .A2(_03626_),
    .ZN(_03632_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07982_ (.A1(_03551_),
    .A2(_03626_),
    .B(_03632_),
    .ZN(_00833_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07983_ (.A1(\u_cpu.rf_ram.memory[116][6] ),
    .A2(_03626_),
    .ZN(_03633_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07984_ (.A1(_03553_),
    .A2(_03626_),
    .B(_03633_),
    .ZN(_00834_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07985_ (.A1(\u_cpu.rf_ram.memory[116][7] ),
    .A2(_03626_),
    .ZN(_03634_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07986_ (.A1(_03555_),
    .A2(_03626_),
    .B(_03634_),
    .ZN(_00835_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07987_ (.A1(_02539_),
    .A2(_02639_),
    .ZN(_03635_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07988_ (.I(_03635_),
    .Z(_03636_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07989_ (.A1(\u_cpu.rf_ram.memory[33][0] ),
    .A2(_03636_),
    .ZN(_03637_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07990_ (.A1(_03539_),
    .A2(_03636_),
    .B(_03637_),
    .ZN(_00836_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07991_ (.A1(\u_cpu.rf_ram.memory[33][1] ),
    .A2(_03636_),
    .ZN(_03638_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07992_ (.A1(_03543_),
    .A2(_03636_),
    .B(_03638_),
    .ZN(_00837_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07993_ (.A1(\u_cpu.rf_ram.memory[33][2] ),
    .A2(_03636_),
    .ZN(_03639_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07994_ (.A1(_03545_),
    .A2(_03636_),
    .B(_03639_),
    .ZN(_00838_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07995_ (.A1(\u_cpu.rf_ram.memory[33][3] ),
    .A2(_03636_),
    .ZN(_03640_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07996_ (.A1(_03547_),
    .A2(_03636_),
    .B(_03640_),
    .ZN(_00839_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07997_ (.A1(\u_cpu.rf_ram.memory[33][4] ),
    .A2(_03636_),
    .ZN(_03641_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07998_ (.A1(_03549_),
    .A2(_03636_),
    .B(_03641_),
    .ZN(_00840_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07999_ (.A1(\u_cpu.rf_ram.memory[33][5] ),
    .A2(_03636_),
    .ZN(_03642_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08000_ (.A1(_03551_),
    .A2(_03636_),
    .B(_03642_),
    .ZN(_00841_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08001_ (.A1(\u_cpu.rf_ram.memory[33][6] ),
    .A2(_03636_),
    .ZN(_03643_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08002_ (.A1(_03553_),
    .A2(_03636_),
    .B(_03643_),
    .ZN(_00842_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08003_ (.A1(\u_cpu.rf_ram.memory[33][7] ),
    .A2(_03636_),
    .ZN(_03644_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08004_ (.A1(_03555_),
    .A2(_03636_),
    .B(_03644_),
    .ZN(_00843_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08005_ (.A1(\u_cpu.cpu.bufreg.lsb[1] ),
    .A2(\u_cpu.cpu.mem_bytecnt[1] ),
    .B(\u_cpu.cpu.mem_bytecnt[0] ),
    .C(\u_cpu.cpu.bufreg.lsb[0] ),
    .ZN(_03645_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08006_ (.A1(\u_cpu.cpu.bufreg.lsb[1] ),
    .A2(\u_cpu.cpu.mem_bytecnt[1] ),
    .ZN(_03646_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08007_ (.A1(_02305_),
    .A2(_03645_),
    .A3(_03646_),
    .ZN(_03647_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08008_ (.A1(_02772_),
    .A2(_03647_),
    .ZN(_03648_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08009_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[0] ),
    .A2(_02774_),
    .ZN(_03649_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08010_ (.A1(_03648_),
    .A2(_03649_),
    .ZN(_03650_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08011_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[1] ),
    .A2(_02774_),
    .B(_02781_),
    .ZN(_03651_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08012_ (.A1(\u_arbiter.i_wb_cpu_ack ),
    .A2(_01442_),
    .Z(_03652_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08013_ (.I(_03652_),
    .Z(_03653_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08014_ (.A1(_03653_),
    .A2(_03648_),
    .ZN(_03654_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08015_ (.A1(\u_arbiter.i_wb_cpu_rdt[0] ),
    .A2(_03653_),
    .B1(_03654_),
    .B2(\u_arbiter.i_wb_cpu_dbus_dat[0] ),
    .ZN(_03655_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08016_ (.A1(_03650_),
    .A2(_03651_),
    .B(_03655_),
    .ZN(_00844_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08017_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[2] ),
    .A2(_02774_),
    .ZN(_03656_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08018_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[0] ),
    .A2(\u_arbiter.i_wb_cpu_dbus_dat[1] ),
    .B(_02774_),
    .ZN(_03657_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08019_ (.A1(_03648_),
    .A2(_03657_),
    .ZN(_03658_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08020_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[1] ),
    .A2(_03650_),
    .ZN(_03659_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08021_ (.A1(_03656_),
    .A2(_03658_),
    .B(_02781_),
    .C(_03659_),
    .ZN(_03660_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08022_ (.A1(\u_arbiter.i_wb_cpu_rdt[1] ),
    .A2(_02781_),
    .B(_03660_),
    .ZN(_03661_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _08023_ (.I(_03661_),
    .ZN(_00845_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08024_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[3] ),
    .A2(_02774_),
    .ZN(_03662_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _08025_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[0] ),
    .A2(\u_arbiter.i_wb_cpu_dbus_dat[1] ),
    .A3(\u_arbiter.i_wb_cpu_dbus_dat[2] ),
    .B(_02774_),
    .ZN(_03663_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08026_ (.A1(_03648_),
    .A2(_03663_),
    .ZN(_03664_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08027_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[2] ),
    .A2(_03658_),
    .ZN(_03665_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08028_ (.A1(_03662_),
    .A2(_03664_),
    .B(_02781_),
    .C(_03665_),
    .ZN(_03666_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08029_ (.A1(\u_arbiter.i_wb_cpu_rdt[2] ),
    .A2(_02781_),
    .B(_03666_),
    .ZN(_03667_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _08030_ (.I(_03667_),
    .ZN(_00846_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08031_ (.I(\u_arbiter.i_wb_cpu_rdt[3] ),
    .ZN(_03668_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08032_ (.I(_03653_),
    .Z(_03669_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08033_ (.A1(_02774_),
    .A2(_02775_),
    .ZN(_03670_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08034_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[4] ),
    .A2(_02774_),
    .B(_03648_),
    .C(_03670_),
    .ZN(_03671_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08035_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[3] ),
    .A2(_03664_),
    .B(_03653_),
    .ZN(_03672_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08036_ (.A1(_03668_),
    .A2(_03669_),
    .B1(_03671_),
    .B2(_03672_),
    .ZN(_00847_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08037_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[4] ),
    .A2(_02775_),
    .Z(_03673_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08038_ (.A1(_02774_),
    .A2(_03673_),
    .ZN(_03674_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08039_ (.A1(_02781_),
    .A2(_03648_),
    .Z(_03675_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08040_ (.I(_03675_),
    .Z(_03676_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08041_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[5] ),
    .A2(_02774_),
    .B(_03674_),
    .C(_03676_),
    .ZN(_03677_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08042_ (.I(_03654_),
    .Z(_03678_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08043_ (.A1(\u_arbiter.i_wb_cpu_rdt[4] ),
    .A2(_03669_),
    .B1(_03678_),
    .B2(\u_arbiter.i_wb_cpu_dbus_dat[4] ),
    .ZN(_03679_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08044_ (.A1(_03677_),
    .A2(_03679_),
    .ZN(_00848_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08045_ (.A1(\u_arbiter.i_wb_cpu_rdt[5] ),
    .A2(_03669_),
    .ZN(_03680_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08046_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[5] ),
    .A2(_03654_),
    .B1(_03676_),
    .B2(_02779_),
    .ZN(_03681_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08047_ (.A1(_03680_),
    .A2(_03681_),
    .ZN(_00849_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _08048_ (.A1(\u_arbiter.i_wb_cpu_rdt[6] ),
    .A2(_03653_),
    .B1(_03654_),
    .B2(\u_arbiter.i_wb_cpu_dbus_dat[6] ),
    .C1(_03676_),
    .C2(\u_arbiter.i_wb_cpu_dbus_dat[7] ),
    .ZN(_03682_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _08049_ (.I(_03682_),
    .ZN(_00850_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08050_ (.I(_03676_),
    .Z(_03683_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08051_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[8] ),
    .A2(_03683_),
    .ZN(_03684_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08052_ (.A1(\u_arbiter.i_wb_cpu_rdt[7] ),
    .A2(_03669_),
    .B1(_03678_),
    .B2(\u_arbiter.i_wb_cpu_dbus_dat[7] ),
    .ZN(_03685_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08053_ (.A1(_03684_),
    .A2(_03685_),
    .ZN(_00851_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08054_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[9] ),
    .A2(_03683_),
    .ZN(_03686_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08055_ (.A1(\u_arbiter.i_wb_cpu_rdt[8] ),
    .A2(_03669_),
    .B1(_03678_),
    .B2(\u_arbiter.i_wb_cpu_dbus_dat[8] ),
    .ZN(_03687_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08056_ (.A1(_03686_),
    .A2(_03687_),
    .ZN(_00852_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08057_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[10] ),
    .A2(_03683_),
    .ZN(_03688_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08058_ (.A1(\u_arbiter.i_wb_cpu_rdt[9] ),
    .A2(_03669_),
    .B1(_03678_),
    .B2(\u_arbiter.i_wb_cpu_dbus_dat[9] ),
    .ZN(_03689_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08059_ (.A1(_03688_),
    .A2(_03689_),
    .ZN(_00853_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08060_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[11] ),
    .A2(_03683_),
    .ZN(_03690_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08061_ (.A1(\u_arbiter.i_wb_cpu_rdt[10] ),
    .A2(_03669_),
    .B1(_03678_),
    .B2(\u_arbiter.i_wb_cpu_dbus_dat[10] ),
    .ZN(_03691_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08062_ (.A1(_03690_),
    .A2(_03691_),
    .ZN(_00854_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08063_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[12] ),
    .A2(_03683_),
    .ZN(_03692_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08064_ (.A1(\u_arbiter.i_wb_cpu_rdt[11] ),
    .A2(_03669_),
    .B1(_03678_),
    .B2(\u_arbiter.i_wb_cpu_dbus_dat[11] ),
    .ZN(_03693_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08065_ (.A1(_03692_),
    .A2(_03693_),
    .ZN(_00855_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08066_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[13] ),
    .A2(_03683_),
    .ZN(_03694_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08067_ (.A1(\u_arbiter.i_wb_cpu_rdt[12] ),
    .A2(_03669_),
    .B1(_03678_),
    .B2(\u_arbiter.i_wb_cpu_dbus_dat[12] ),
    .ZN(_03695_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08068_ (.A1(_03694_),
    .A2(_03695_),
    .ZN(_00856_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08069_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[14] ),
    .A2(_03683_),
    .ZN(_03696_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08070_ (.A1(\u_arbiter.i_wb_cpu_rdt[13] ),
    .A2(_03669_),
    .B1(_03678_),
    .B2(\u_arbiter.i_wb_cpu_dbus_dat[13] ),
    .ZN(_03697_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08071_ (.A1(_03696_),
    .A2(_03697_),
    .ZN(_00857_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _08072_ (.A1(\u_arbiter.i_wb_cpu_rdt[14] ),
    .A2(_03653_),
    .B1(_03654_),
    .B2(\u_arbiter.i_wb_cpu_dbus_dat[14] ),
    .C1(_03676_),
    .C2(\u_arbiter.i_wb_cpu_dbus_dat[15] ),
    .ZN(_03698_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _08073_ (.I(_03698_),
    .ZN(_00858_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08074_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[16] ),
    .A2(_03683_),
    .ZN(_03699_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08075_ (.A1(\u_arbiter.i_wb_cpu_rdt[15] ),
    .A2(_03669_),
    .B1(_03678_),
    .B2(\u_arbiter.i_wb_cpu_dbus_dat[15] ),
    .ZN(_03700_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08076_ (.A1(_03699_),
    .A2(_03700_),
    .ZN(_00859_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08077_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[17] ),
    .A2(_03683_),
    .ZN(_03701_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08078_ (.A1(\u_arbiter.i_wb_cpu_rdt[16] ),
    .A2(_03669_),
    .B1(_03678_),
    .B2(\u_arbiter.i_wb_cpu_dbus_dat[16] ),
    .ZN(_03702_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08079_ (.A1(_03701_),
    .A2(_03702_),
    .ZN(_00860_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _08080_ (.A1(\u_arbiter.i_wb_cpu_rdt[17] ),
    .A2(_03653_),
    .B1(_03654_),
    .B2(\u_arbiter.i_wb_cpu_dbus_dat[17] ),
    .C1(_03676_),
    .C2(\u_arbiter.i_wb_cpu_dbus_dat[18] ),
    .ZN(_03703_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _08081_ (.I(_03703_),
    .ZN(_00861_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08082_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[19] ),
    .A2(_03683_),
    .ZN(_03704_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08083_ (.A1(\u_arbiter.i_wb_cpu_rdt[18] ),
    .A2(_03669_),
    .B1(_03678_),
    .B2(\u_arbiter.i_wb_cpu_dbus_dat[18] ),
    .ZN(_03705_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08084_ (.A1(_03704_),
    .A2(_03705_),
    .ZN(_00862_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08085_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[20] ),
    .A2(_03683_),
    .ZN(_03706_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08086_ (.A1(\u_arbiter.i_wb_cpu_rdt[19] ),
    .A2(_03669_),
    .B1(_03678_),
    .B2(\u_arbiter.i_wb_cpu_dbus_dat[19] ),
    .ZN(_03707_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08087_ (.A1(_03706_),
    .A2(_03707_),
    .ZN(_00863_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08088_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[21] ),
    .A2(_03683_),
    .ZN(_03708_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08089_ (.A1(\u_arbiter.i_wb_cpu_rdt[20] ),
    .A2(_03669_),
    .B1(_03654_),
    .B2(\u_arbiter.i_wb_cpu_dbus_dat[20] ),
    .ZN(_03709_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08090_ (.A1(_03708_),
    .A2(_03709_),
    .ZN(_00864_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _08091_ (.A1(\u_arbiter.i_wb_cpu_rdt[21] ),
    .A2(_03653_),
    .B1(_03654_),
    .B2(\u_arbiter.i_wb_cpu_dbus_dat[21] ),
    .C1(_03676_),
    .C2(\u_arbiter.i_wb_cpu_dbus_dat[22] ),
    .ZN(_03710_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _08092_ (.I(_03710_),
    .ZN(_00865_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08093_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[23] ),
    .A2(_03683_),
    .ZN(_03711_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08094_ (.A1(\u_arbiter.i_wb_cpu_rdt[22] ),
    .A2(_03653_),
    .B1(_03654_),
    .B2(\u_arbiter.i_wb_cpu_dbus_dat[22] ),
    .ZN(_03712_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08095_ (.A1(_03711_),
    .A2(_03712_),
    .ZN(_00866_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08096_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[24] ),
    .A2(_03683_),
    .ZN(_03713_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08097_ (.A1(\u_arbiter.i_wb_cpu_rdt[23] ),
    .A2(_03653_),
    .B1(_03654_),
    .B2(\u_arbiter.i_wb_cpu_dbus_dat[23] ),
    .ZN(_03714_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08098_ (.A1(_03713_),
    .A2(_03714_),
    .ZN(_00867_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08099_ (.A1(\u_arbiter.i_wb_cpu_rdt[24] ),
    .A2(_03669_),
    .ZN(_03715_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08100_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[24] ),
    .A2(_03654_),
    .B1(_03676_),
    .B2(\u_arbiter.i_wb_cpu_dbus_dat[25] ),
    .ZN(_03716_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08101_ (.A1(_03715_),
    .A2(_03716_),
    .ZN(_00868_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08102_ (.I(\u_arbiter.i_wb_cpu_dbus_dat[26] ),
    .ZN(_03717_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08103_ (.A1(_02781_),
    .A2(_03648_),
    .ZN(_03718_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08104_ (.A1(\u_arbiter.i_wb_cpu_rdt[25] ),
    .A2(_03653_),
    .B1(_03654_),
    .B2(\u_arbiter.i_wb_cpu_dbus_dat[25] ),
    .ZN(_03719_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08105_ (.A1(_03717_),
    .A2(_03718_),
    .B(_03719_),
    .ZN(_00869_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _08106_ (.A1(\u_arbiter.i_wb_cpu_rdt[26] ),
    .A2(_02781_),
    .B1(_03718_),
    .B2(\u_arbiter.i_wb_cpu_dbus_dat[27] ),
    .ZN(_03720_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08107_ (.A1(_03717_),
    .A2(_03678_),
    .B(_03720_),
    .ZN(_00870_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08108_ (.A1(\u_arbiter.i_wb_cpu_dbus_dat[28] ),
    .A2(_03676_),
    .ZN(_03721_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08109_ (.A1(\u_arbiter.i_wb_cpu_rdt[27] ),
    .A2(_03653_),
    .B1(_03654_),
    .B2(\u_arbiter.i_wb_cpu_dbus_dat[27] ),
    .ZN(_03722_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08110_ (.A1(_03721_),
    .A2(_03722_),
    .ZN(_00871_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08111_ (.I(\u_arbiter.i_wb_cpu_dbus_dat[29] ),
    .ZN(_03723_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08112_ (.A1(\u_arbiter.i_wb_cpu_rdt[28] ),
    .A2(_03653_),
    .B1(_03654_),
    .B2(\u_arbiter.i_wb_cpu_dbus_dat[28] ),
    .ZN(_03724_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08113_ (.A1(_03723_),
    .A2(_03718_),
    .B(_03724_),
    .ZN(_00872_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08114_ (.I(\u_arbiter.i_wb_cpu_dbus_dat[30] ),
    .ZN(_03725_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08115_ (.A1(\u_arbiter.i_wb_cpu_rdt[29] ),
    .A2(_02781_),
    .ZN(_03726_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _08116_ (.A1(_03723_),
    .A2(_03678_),
    .B1(_03683_),
    .B2(_03725_),
    .C(_03726_),
    .ZN(_00873_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08117_ (.I(\u_arbiter.i_wb_cpu_dbus_dat[31] ),
    .ZN(_03727_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08118_ (.A1(\u_arbiter.i_wb_cpu_rdt[30] ),
    .A2(_02781_),
    .ZN(_03728_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _08119_ (.A1(_03725_),
    .A2(_03678_),
    .B1(_03683_),
    .B2(_03727_),
    .C(_03728_),
    .ZN(_00874_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _08120_ (.A1(\u_arbiter.i_wb_cpu_rdt[31] ),
    .A2(_02781_),
    .B1(_03718_),
    .B2(_02325_),
    .ZN(_03729_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08121_ (.A1(_03727_),
    .A2(_03678_),
    .B(_03729_),
    .ZN(_00875_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08122_ (.A1(_02539_),
    .A2(_02821_),
    .ZN(_03730_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08123_ (.I(_03730_),
    .Z(_03731_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08124_ (.A1(\u_cpu.rf_ram.memory[113][0] ),
    .A2(_03731_),
    .ZN(_03732_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08125_ (.A1(_03539_),
    .A2(_03731_),
    .B(_03732_),
    .ZN(_00876_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08126_ (.A1(\u_cpu.rf_ram.memory[113][1] ),
    .A2(_03731_),
    .ZN(_03733_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08127_ (.A1(_03543_),
    .A2(_03731_),
    .B(_03733_),
    .ZN(_00877_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08128_ (.A1(\u_cpu.rf_ram.memory[113][2] ),
    .A2(_03731_),
    .ZN(_03734_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08129_ (.A1(_03545_),
    .A2(_03731_),
    .B(_03734_),
    .ZN(_00878_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08130_ (.A1(\u_cpu.rf_ram.memory[113][3] ),
    .A2(_03731_),
    .ZN(_03735_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08131_ (.A1(_03547_),
    .A2(_03731_),
    .B(_03735_),
    .ZN(_00879_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08132_ (.A1(\u_cpu.rf_ram.memory[113][4] ),
    .A2(_03731_),
    .ZN(_03736_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08133_ (.A1(_03549_),
    .A2(_03731_),
    .B(_03736_),
    .ZN(_00880_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08134_ (.A1(\u_cpu.rf_ram.memory[113][5] ),
    .A2(_03731_),
    .ZN(_03737_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08135_ (.A1(_03551_),
    .A2(_03731_),
    .B(_03737_),
    .ZN(_00881_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08136_ (.A1(\u_cpu.rf_ram.memory[113][6] ),
    .A2(_03731_),
    .ZN(_03738_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08137_ (.A1(_03553_),
    .A2(_03731_),
    .B(_03738_),
    .ZN(_00882_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08138_ (.A1(\u_cpu.rf_ram.memory[113][7] ),
    .A2(_03731_),
    .ZN(_03739_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08139_ (.A1(_03555_),
    .A2(_03731_),
    .B(_03739_),
    .ZN(_00883_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08140_ (.I(_02768_),
    .Z(_03740_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08141_ (.I0(\u_arbiter.i_wb_cpu_rdt[11] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[11] ),
    .S(_01434_),
    .Z(_03741_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08142_ (.I0(\u_arbiter.i_wb_cpu_rdt[10] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[10] ),
    .S(_01434_),
    .Z(_03742_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08143_ (.I0(\u_arbiter.i_wb_cpu_rdt[9] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[9] ),
    .S(_01435_),
    .Z(_03743_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08144_ (.I0(\u_arbiter.i_wb_cpu_rdt[7] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[7] ),
    .S(_01434_),
    .Z(_03744_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _08145_ (.A1(_03741_),
    .A2(_03742_),
    .A3(_03743_),
    .A4(_03744_),
    .ZN(_03745_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08146_ (.A1(_01436_),
    .A2(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[8] ),
    .Z(_03746_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08147_ (.A1(_02765_),
    .A2(\u_arbiter.i_wb_cpu_rdt[8] ),
    .B(_03746_),
    .ZN(_03747_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08148_ (.A1(_03745_),
    .A2(_03747_),
    .Z(_03748_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08149_ (.I(_03748_),
    .ZN(_03749_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08150_ (.A1(_01436_),
    .A2(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[12] ),
    .Z(_03750_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08151_ (.A1(_02765_),
    .A2(\u_arbiter.i_wb_cpu_rdt[12] ),
    .B(_03750_),
    .ZN(_03751_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08152_ (.A1(_03749_),
    .A2(_03751_),
    .ZN(_03752_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08153_ (.A1(_01436_),
    .A2(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[0] ),
    .Z(_03753_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08154_ (.A1(_02765_),
    .A2(\u_arbiter.i_wb_cpu_rdt[0] ),
    .B(_03753_),
    .ZN(_03754_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08155_ (.I0(\u_arbiter.i_wb_cpu_rdt[1] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[1] ),
    .S(_01435_),
    .Z(_03755_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08156_ (.I0(\u_arbiter.i_wb_cpu_rdt[6] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[6] ),
    .S(_01435_),
    .Z(_03756_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08157_ (.I(_03756_),
    .ZN(_03757_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08158_ (.A1(_01436_),
    .A2(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[5] ),
    .Z(_03758_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08159_ (.A1(_02765_),
    .A2(\u_arbiter.i_wb_cpu_rdt[5] ),
    .B(_03758_),
    .ZN(_03759_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08160_ (.A1(_01435_),
    .A2(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[3] ),
    .ZN(_03760_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08161_ (.A1(_01435_),
    .A2(_03668_),
    .B(_03760_),
    .ZN(_03761_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08162_ (.I0(\u_arbiter.i_wb_cpu_rdt[4] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[4] ),
    .S(_01435_),
    .Z(_03762_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08163_ (.I0(\u_arbiter.i_wb_cpu_rdt[2] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[2] ),
    .S(_01435_),
    .Z(_03763_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _08164_ (.A1(_03761_),
    .A2(_03762_),
    .A3(_03763_),
    .ZN(_03764_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08165_ (.A1(_03757_),
    .A2(_03759_),
    .A3(_03764_),
    .ZN(_03765_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08166_ (.A1(_01435_),
    .A2(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[14] ),
    .Z(_03766_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08167_ (.A1(_02765_),
    .A2(\u_arbiter.i_wb_cpu_rdt[14] ),
    .B(_03766_),
    .ZN(_03767_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08168_ (.I0(\u_arbiter.i_wb_cpu_rdt[15] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[15] ),
    .S(_01436_),
    .Z(_03768_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08169_ (.A1(_03767_),
    .A2(_03768_),
    .ZN(_03769_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08170_ (.A1(_03765_),
    .A2(_03769_),
    .ZN(_03770_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08171_ (.A1(_03754_),
    .A2(_03755_),
    .A3(_03770_),
    .ZN(_03771_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08172_ (.I0(\u_arbiter.i_wb_cpu_rdt[0] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[0] ),
    .S(_01435_),
    .Z(_03772_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08173_ (.I(_03772_),
    .Z(_03773_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08174_ (.A1(_03773_),
    .A2(_03755_),
    .ZN(_03774_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08175_ (.I0(\u_arbiter.i_wb_cpu_rdt[14] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[14] ),
    .S(_01435_),
    .Z(_03775_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08176_ (.I(_03775_),
    .Z(_03776_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08177_ (.A1(_01435_),
    .A2(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[15] ),
    .Z(_03777_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08178_ (.A1(_02765_),
    .A2(\u_arbiter.i_wb_cpu_rdt[15] ),
    .B(_03777_),
    .ZN(_03778_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08179_ (.A1(_03776_),
    .A2(_03778_),
    .ZN(_03779_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08180_ (.A1(_03773_),
    .A2(_03755_),
    .ZN(_03780_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08181_ (.A1(_03779_),
    .A2(_03780_),
    .ZN(_03781_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08182_ (.A1(_03774_),
    .A2(_03781_),
    .ZN(_03782_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08183_ (.A1(_03763_),
    .A2(_03782_),
    .ZN(_03783_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08184_ (.A1(_01435_),
    .A2(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[13] ),
    .Z(_03784_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08185_ (.A1(_02765_),
    .A2(\u_arbiter.i_wb_cpu_rdt[13] ),
    .B(_03784_),
    .ZN(_03785_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08186_ (.A1(_03776_),
    .A2(_03785_),
    .ZN(_03786_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08187_ (.A1(_03776_),
    .A2(_03778_),
    .ZN(_03787_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08188_ (.I0(\u_arbiter.i_wb_cpu_rdt[8] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[8] ),
    .S(_01435_),
    .Z(_03788_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08189_ (.A1(_03745_),
    .A2(_03788_),
    .Z(_03789_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _08190_ (.A1(_03785_),
    .A2(_03787_),
    .A3(_03789_),
    .ZN(_03790_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08191_ (.A1(_03754_),
    .A2(_03755_),
    .ZN(_03791_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08192_ (.A1(_03786_),
    .A2(_03790_),
    .B(_03791_),
    .ZN(_03792_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08193_ (.A1(_03752_),
    .A2(_03771_),
    .B(_03783_),
    .C(_03792_),
    .ZN(_03793_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08194_ (.A1(_03740_),
    .A2(_03793_),
    .ZN(_03794_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08195_ (.A1(_02383_),
    .A2(_03740_),
    .B(_03794_),
    .ZN(_00884_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08196_ (.A1(_02765_),
    .A2(\u_arbiter.i_wb_cpu_ibus_adr[1] ),
    .ZN(_03795_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08197_ (.A1(\u_arbiter.i_wb_cpu_ack ),
    .A2(_01431_),
    .A3(_03795_),
    .ZN(_03796_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08198_ (.I(_03796_),
    .Z(_03797_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08199_ (.I(_03797_),
    .Z(_03798_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08200_ (.A1(_01436_),
    .A2(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[1] ),
    .Z(_03799_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08201_ (.A1(_02765_),
    .A2(\u_arbiter.i_wb_cpu_rdt[1] ),
    .B(_03799_),
    .ZN(_03800_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08202_ (.A1(_03773_),
    .A2(_03800_),
    .ZN(_03801_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08203_ (.I0(\u_arbiter.i_wb_cpu_rdt[13] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[13] ),
    .S(_01436_),
    .Z(_03802_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08204_ (.A1(_03767_),
    .A2(_03802_),
    .ZN(_03803_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08205_ (.A1(_03801_),
    .A2(_03803_),
    .ZN(_03804_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08206_ (.A1(_03761_),
    .A2(_03782_),
    .B(_03804_),
    .ZN(_03805_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08207_ (.A1(\u_cpu.cpu.decode.opcode[1] ),
    .A2(_03798_),
    .ZN(_03806_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08208_ (.A1(_03798_),
    .A2(_03805_),
    .B(_03806_),
    .ZN(_00885_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _08209_ (.A1(_03765_),
    .A2(_03778_),
    .Z(_03807_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _08210_ (.A1(_03752_),
    .A2(_03800_),
    .A3(_03807_),
    .Z(_03808_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08211_ (.A1(_03776_),
    .A2(_03768_),
    .ZN(_03809_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08212_ (.A1(_03803_),
    .A2(_03809_),
    .ZN(_03810_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08213_ (.A1(_03774_),
    .A2(_03781_),
    .Z(_03811_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08214_ (.A1(_02768_),
    .A2(_03811_),
    .ZN(_03812_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08215_ (.A1(_03773_),
    .A2(_03810_),
    .B(_03812_),
    .ZN(_03813_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08216_ (.A1(_03773_),
    .A2(_03767_),
    .B(_03808_),
    .C(_03813_),
    .ZN(_03814_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08217_ (.A1(_03796_),
    .A2(_03811_),
    .ZN(_03815_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08218_ (.I(_03815_),
    .Z(_03816_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08219_ (.A1(_01372_),
    .A2(_03798_),
    .B1(_03762_),
    .B2(_03816_),
    .ZN(_03817_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08220_ (.A1(_03814_),
    .A2(_03817_),
    .ZN(_00886_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08221_ (.A1(_03769_),
    .A2(_03802_),
    .ZN(_03818_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08222_ (.A1(_03741_),
    .A2(_03742_),
    .Z(_03819_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08223_ (.A1(_03818_),
    .A2(_03819_),
    .B(_03790_),
    .C(_03810_),
    .ZN(_03820_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08224_ (.A1(_03791_),
    .A2(_03820_),
    .ZN(_03821_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _08225_ (.A1(_03754_),
    .A2(_03778_),
    .B1(_03782_),
    .B2(_03759_),
    .C(_03797_),
    .ZN(_03822_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08226_ (.A1(_02306_),
    .A2(_03798_),
    .B1(_03821_),
    .B2(_03822_),
    .ZN(_03823_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _08227_ (.I(_03823_),
    .ZN(_00887_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08228_ (.A1(_01374_),
    .A2(_02768_),
    .ZN(_03824_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _08229_ (.A1(_03771_),
    .A2(_03813_),
    .B1(_03816_),
    .B2(_03757_),
    .C(_03824_),
    .ZN(_00888_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08230_ (.A1(_03754_),
    .A2(_03755_),
    .ZN(_03825_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08231_ (.A1(_03767_),
    .A2(_03778_),
    .ZN(_03826_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08232_ (.A1(_03757_),
    .A2(_03759_),
    .B(_03819_),
    .ZN(_03827_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08233_ (.A1(_03767_),
    .A2(_03778_),
    .ZN(_03828_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _08234_ (.A1(_03763_),
    .A2(_03790_),
    .B1(_03818_),
    .B2(_03827_),
    .C1(_03828_),
    .C2(_03802_),
    .ZN(_03829_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08235_ (.I0(\u_arbiter.i_wb_cpu_rdt[12] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[12] ),
    .S(_01435_),
    .Z(_03830_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08236_ (.I(_03830_),
    .Z(_03831_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08237_ (.A1(_03782_),
    .A2(_03804_),
    .B(_03831_),
    .ZN(_03832_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _08238_ (.A1(_03825_),
    .A2(_03826_),
    .B1(_03829_),
    .B2(_03801_),
    .C(_03832_),
    .ZN(_03833_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08239_ (.A1(_03740_),
    .A2(_03833_),
    .ZN(_03834_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08240_ (.A1(_02333_),
    .A2(_03740_),
    .B(_03834_),
    .ZN(_00889_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08241_ (.A1(_03751_),
    .A2(_03803_),
    .ZN(_03835_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08242_ (.A1(_03741_),
    .A2(_03818_),
    .ZN(_03836_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08243_ (.A1(_03742_),
    .A2(_03757_),
    .B(_03836_),
    .ZN(_03837_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08244_ (.A1(_03761_),
    .A2(_03790_),
    .B(_03835_),
    .C(_03837_),
    .ZN(_03838_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _08245_ (.A1(_03773_),
    .A2(_03767_),
    .B1(_03801_),
    .B2(_03838_),
    .C(_03811_),
    .ZN(_03839_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08246_ (.A1(_03811_),
    .A2(_03802_),
    .B(_03839_),
    .C(_02768_),
    .ZN(_03840_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08247_ (.A1(_02332_),
    .A2(_03740_),
    .B(_03840_),
    .ZN(_00890_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _08248_ (.A1(_03757_),
    .A2(_03759_),
    .A3(_03819_),
    .Z(_03841_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08249_ (.I(_03841_),
    .ZN(_03842_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _08250_ (.A1(_03762_),
    .A2(_03790_),
    .B1(_03818_),
    .B2(_03842_),
    .C(_03835_),
    .ZN(_03843_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _08251_ (.A1(_03767_),
    .A2(_03774_),
    .B1(_03801_),
    .B2(_03843_),
    .ZN(_03844_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08252_ (.A1(_03740_),
    .A2(_03844_),
    .ZN(_03845_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08253_ (.A1(_01408_),
    .A2(_03740_),
    .B(_03845_),
    .ZN(_00891_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08254_ (.I0(\u_arbiter.i_wb_cpu_rdt[20] ),
    .I1(\u_arbiter.i_wb_cpu_rdt[4] ),
    .S(_01437_),
    .Z(_03846_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _08255_ (.A1(_03752_),
    .A2(_03770_),
    .B1(_03787_),
    .B2(_03763_),
    .C(_03800_),
    .ZN(_03847_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08256_ (.A1(_03763_),
    .A2(_03785_),
    .A3(_03809_),
    .ZN(_03848_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08257_ (.A1(_03786_),
    .A2(_03790_),
    .B(_03831_),
    .ZN(_03849_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _08258_ (.A1(_03773_),
    .A2(_03848_),
    .A3(_03849_),
    .Z(_03850_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08259_ (.A1(_03754_),
    .A2(_03800_),
    .ZN(_03851_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08260_ (.A1(_03763_),
    .A2(_03828_),
    .B(_03851_),
    .ZN(_03852_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08261_ (.A1(_02768_),
    .A2(_03774_),
    .ZN(_03853_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _08262_ (.A1(_03847_),
    .A2(_03850_),
    .A3(_03852_),
    .A4(_03853_),
    .ZN(_03854_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08263_ (.A1(_03816_),
    .A2(_03846_),
    .B(_03854_),
    .ZN(_03855_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08264_ (.A1(_01381_),
    .A2(_03740_),
    .B(_03855_),
    .ZN(_00892_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08265_ (.I0(\u_arbiter.i_wb_cpu_rdt[21] ),
    .I1(\u_arbiter.i_wb_cpu_rdt[5] ),
    .S(_01437_),
    .Z(_03856_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08266_ (.A1(_03761_),
    .A2(_03828_),
    .ZN(_03857_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08267_ (.A1(_03831_),
    .A2(_03790_),
    .ZN(_03858_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08268_ (.A1(_03773_),
    .A2(_03858_),
    .ZN(_03859_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08269_ (.A1(_03767_),
    .A2(_03768_),
    .ZN(_03860_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08270_ (.A1(_03768_),
    .A2(_03802_),
    .ZN(_03861_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08271_ (.A1(_03767_),
    .A2(_03861_),
    .ZN(_03862_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _08272_ (.A1(_03773_),
    .A2(_03860_),
    .B1(_03862_),
    .B2(_03755_),
    .ZN(_03863_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08273_ (.A1(_03800_),
    .A2(_03859_),
    .B1(_03863_),
    .B2(_03761_),
    .ZN(_03864_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08274_ (.A1(_03780_),
    .A2(_03857_),
    .B(_03864_),
    .ZN(_03865_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08275_ (.A1(_03816_),
    .A2(_03856_),
    .B1(_03865_),
    .B2(_02768_),
    .ZN(_03866_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08276_ (.A1(_02343_),
    .A2(_03740_),
    .B(_03866_),
    .ZN(_00893_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08277_ (.I0(\u_arbiter.i_wb_cpu_rdt[22] ),
    .I1(\u_arbiter.i_wb_cpu_rdt[6] ),
    .S(_01436_),
    .Z(_03867_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08278_ (.A1(_03801_),
    .A2(_03858_),
    .ZN(_03868_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08279_ (.A1(_03858_),
    .A2(_03862_),
    .ZN(_03869_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08280_ (.A1(_03791_),
    .A2(_03869_),
    .ZN(_03870_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08281_ (.A1(_03825_),
    .A2(_03870_),
    .ZN(_03871_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08282_ (.A1(_03762_),
    .A2(_03868_),
    .B(_03871_),
    .ZN(_03872_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08283_ (.A1(_03762_),
    .A2(_03828_),
    .ZN(_03873_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _08284_ (.A1(_03756_),
    .A2(_03778_),
    .B1(_03779_),
    .B2(_03867_),
    .C(_03851_),
    .ZN(_03874_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08285_ (.A1(_03851_),
    .A2(_03872_),
    .B1(_03873_),
    .B2(_03874_),
    .ZN(_03875_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08286_ (.A1(_03796_),
    .A2(_03782_),
    .ZN(_03876_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08287_ (.A1(_03816_),
    .A2(_03867_),
    .B1(_03875_),
    .B2(_03876_),
    .ZN(_03877_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08288_ (.A1(_02337_),
    .A2(_03740_),
    .B(_03877_),
    .ZN(_00894_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08289_ (.A1(_02469_),
    .A2(_02821_),
    .ZN(_03878_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08290_ (.I(_03878_),
    .Z(_03879_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08291_ (.A1(\u_cpu.rf_ram.memory[114][0] ),
    .A2(_03879_),
    .ZN(_03880_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08292_ (.A1(_03539_),
    .A2(_03879_),
    .B(_03880_),
    .ZN(_00895_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08293_ (.A1(\u_cpu.rf_ram.memory[114][1] ),
    .A2(_03879_),
    .ZN(_03881_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08294_ (.A1(_03543_),
    .A2(_03879_),
    .B(_03881_),
    .ZN(_00896_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08295_ (.A1(\u_cpu.rf_ram.memory[114][2] ),
    .A2(_03879_),
    .ZN(_03882_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08296_ (.A1(_03545_),
    .A2(_03879_),
    .B(_03882_),
    .ZN(_00897_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08297_ (.A1(\u_cpu.rf_ram.memory[114][3] ),
    .A2(_03879_),
    .ZN(_03883_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08298_ (.A1(_03547_),
    .A2(_03879_),
    .B(_03883_),
    .ZN(_00898_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08299_ (.A1(\u_cpu.rf_ram.memory[114][4] ),
    .A2(_03879_),
    .ZN(_03884_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08300_ (.A1(_03549_),
    .A2(_03879_),
    .B(_03884_),
    .ZN(_00899_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08301_ (.A1(\u_cpu.rf_ram.memory[114][5] ),
    .A2(_03879_),
    .ZN(_03885_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08302_ (.A1(_03551_),
    .A2(_03879_),
    .B(_03885_),
    .ZN(_00900_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08303_ (.A1(\u_cpu.rf_ram.memory[114][6] ),
    .A2(_03879_),
    .ZN(_03886_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08304_ (.A1(_03553_),
    .A2(_03879_),
    .B(_03886_),
    .ZN(_00901_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08305_ (.A1(\u_cpu.rf_ram.memory[114][7] ),
    .A2(_03879_),
    .ZN(_03887_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08306_ (.A1(_03555_),
    .A2(_03879_),
    .B(_03887_),
    .ZN(_00902_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08307_ (.I0(\u_arbiter.i_wb_cpu_rdt[26] ),
    .I1(\u_arbiter.i_wb_cpu_rdt[10] ),
    .S(_01436_),
    .Z(_03888_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08308_ (.A1(_03816_),
    .A2(_03888_),
    .ZN(_03889_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08309_ (.I0(\u_arbiter.i_wb_cpu_rdt[5] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[5] ),
    .S(_01436_),
    .Z(_03890_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08310_ (.A1(_03745_),
    .A2(_03788_),
    .ZN(_03891_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08311_ (.A1(_03785_),
    .A2(_03787_),
    .ZN(_03892_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08312_ (.A1(_03831_),
    .A2(_03789_),
    .B(_03892_),
    .ZN(_03893_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08313_ (.I(_03893_),
    .ZN(_03894_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08314_ (.A1(_03890_),
    .A2(_03891_),
    .B(_03894_),
    .ZN(_03895_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08315_ (.A1(_03776_),
    .A2(_03768_),
    .ZN(_03896_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08316_ (.A1(_03785_),
    .A2(_03896_),
    .ZN(_03897_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08317_ (.A1(_03831_),
    .A2(_03776_),
    .ZN(_03898_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08318_ (.I(_03898_),
    .ZN(_03899_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08319_ (.A1(_03779_),
    .A2(_03785_),
    .ZN(_03900_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08320_ (.A1(_03741_),
    .A2(_03831_),
    .ZN(_03901_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _08321_ (.A1(_03742_),
    .A2(_03900_),
    .A3(_03901_),
    .ZN(_03902_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08322_ (.A1(_03861_),
    .A2(_03899_),
    .B(_03902_),
    .ZN(_03903_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08323_ (.A1(_03897_),
    .A2(_03903_),
    .ZN(_03904_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _08324_ (.A1(_03744_),
    .A2(_03786_),
    .B1(_03828_),
    .B2(_03890_),
    .C(_03904_),
    .ZN(_03905_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08325_ (.A1(_03831_),
    .A2(_03897_),
    .B(_03791_),
    .ZN(_03906_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08326_ (.A1(_03895_),
    .A2(_03905_),
    .B(_03906_),
    .ZN(_03907_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _08327_ (.A1(_03763_),
    .A2(_03860_),
    .B1(_03828_),
    .B2(_03744_),
    .C(_03800_),
    .ZN(_03908_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08328_ (.A1(_03773_),
    .A2(_03908_),
    .ZN(_03909_));
 gf180mcu_fd_sc_mcu7t5v0__oai222_1 _08329_ (.A1(_03767_),
    .A2(_03890_),
    .B1(_03769_),
    .B2(_03888_),
    .C1(_03826_),
    .C2(_03744_),
    .ZN(_03910_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08330_ (.A1(_03780_),
    .A2(_03910_),
    .ZN(_03911_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08331_ (.A1(_03907_),
    .A2(_03909_),
    .B(_03911_),
    .C(_03876_),
    .ZN(_03912_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08332_ (.A1(_03889_),
    .A2(_03912_),
    .Z(_03913_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08333_ (.A1(_01380_),
    .A2(_03740_),
    .B(_03913_),
    .ZN(_00903_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _08334_ (.A1(_02436_),
    .A2(_02313_),
    .A3(_01376_),
    .B(_02305_),
    .ZN(_03914_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08335_ (.A1(_03796_),
    .A2(_03914_),
    .Z(_03915_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08336_ (.I(_03915_),
    .Z(_03916_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08337_ (.A1(\u_cpu.cpu.immdec.imm24_20[1] ),
    .A2(_03798_),
    .ZN(_03917_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08338_ (.A1(\u_cpu.cpu.immdec.imm24_20[0] ),
    .A2(_03916_),
    .ZN(_03918_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08339_ (.A1(_03916_),
    .A2(_03917_),
    .B(_03918_),
    .C(_03855_),
    .ZN(_00904_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08340_ (.A1(_02768_),
    .A2(_03914_),
    .ZN(_03919_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08341_ (.A1(\u_cpu.cpu.immdec.imm24_20[1] ),
    .A2(_03916_),
    .B1(_03919_),
    .B2(\u_cpu.cpu.immdec.imm24_20[2] ),
    .ZN(_03920_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08342_ (.A1(_03866_),
    .A2(_03920_),
    .ZN(_00905_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08343_ (.I(\u_cpu.cpu.immdec.imm24_20[2] ),
    .ZN(_03921_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08344_ (.A1(\u_cpu.cpu.immdec.imm24_20[3] ),
    .A2(_03914_),
    .B(_03797_),
    .ZN(_03922_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08345_ (.A1(_03921_),
    .A2(_03916_),
    .B1(_03922_),
    .B2(_03877_),
    .ZN(_00906_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08346_ (.I0(\u_arbiter.i_wb_cpu_rdt[23] ),
    .I1(\u_arbiter.i_wb_cpu_rdt[7] ),
    .S(_01436_),
    .Z(_03923_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08347_ (.A1(_03831_),
    .A2(_03790_),
    .B1(_03818_),
    .B2(_03819_),
    .ZN(_03924_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08348_ (.A1(_03870_),
    .A2(_03924_),
    .B(_03759_),
    .ZN(_03925_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08349_ (.A1(_03871_),
    .A2(_03925_),
    .ZN(_03926_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _08350_ (.A1(_03742_),
    .A2(_03768_),
    .Z(_03927_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08351_ (.A1(_03776_),
    .A2(_03923_),
    .B(_03927_),
    .C(_03826_),
    .ZN(_03928_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08352_ (.A1(_03890_),
    .A2(_03896_),
    .B(_03851_),
    .ZN(_03929_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _08353_ (.A1(_03851_),
    .A2(_03926_),
    .B1(_03928_),
    .B2(_03929_),
    .C(_03782_),
    .ZN(_03930_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08354_ (.A1(_03782_),
    .A2(_03923_),
    .B(_03930_),
    .C(_03797_),
    .ZN(_03931_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08355_ (.A1(\u_cpu.cpu.immdec.imm24_20[4] ),
    .A2(_02768_),
    .ZN(_03932_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08356_ (.A1(\u_cpu.cpu.immdec.imm24_20[3] ),
    .A2(_03916_),
    .ZN(_03933_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _08357_ (.A1(_03916_),
    .A2(_03931_),
    .A3(_03932_),
    .B(_03933_),
    .ZN(_00907_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _08358_ (.A1(_03741_),
    .A2(_03786_),
    .B1(_03820_),
    .B2(_03756_),
    .C(_03859_),
    .ZN(_03934_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08359_ (.I0(\u_arbiter.i_wb_cpu_rdt[24] ),
    .I1(\u_arbiter.i_wb_cpu_rdt[8] ),
    .S(_01437_),
    .Z(_03935_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08360_ (.A1(_03741_),
    .A2(_03778_),
    .B1(_03779_),
    .B2(_03935_),
    .ZN(_03936_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08361_ (.A1(_03755_),
    .A2(_03757_),
    .B1(_03780_),
    .B2(_03936_),
    .ZN(_03937_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08362_ (.A1(_03876_),
    .A2(_03937_),
    .ZN(_03938_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _08363_ (.A1(\u_cpu.cpu.immdec.imm24_20[4] ),
    .A2(_03916_),
    .B1(_03919_),
    .B2(\u_cpu.cpu.immdec.imm30_25[0] ),
    .C1(_03935_),
    .C2(_03816_),
    .ZN(_03939_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08364_ (.A1(_03934_),
    .A2(_03938_),
    .B(_03939_),
    .ZN(_00908_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08365_ (.A1(_03773_),
    .A2(_03767_),
    .ZN(_03940_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08366_ (.A1(_03785_),
    .A2(_03891_),
    .ZN(_03941_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08367_ (.A1(_03810_),
    .A2(_03941_),
    .B(_03763_),
    .ZN(_03942_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08368_ (.A1(_03831_),
    .A2(_03861_),
    .B(_03902_),
    .ZN(_03943_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _08369_ (.A1(_03773_),
    .A2(_03858_),
    .A3(_03942_),
    .A4(_03943_),
    .ZN(_03944_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _08370_ (.A1(_03831_),
    .A2(_03773_),
    .B1(_03800_),
    .B2(_03940_),
    .C(_03944_),
    .ZN(_03945_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08371_ (.A1(_03876_),
    .A2(_03945_),
    .Z(_03946_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08372_ (.A1(_02436_),
    .A2(_02313_),
    .A3(_02434_),
    .ZN(_03947_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08373_ (.A1(_02305_),
    .A2(_03947_),
    .ZN(_03948_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08374_ (.A1(_03797_),
    .A2(_03948_),
    .ZN(_03949_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08375_ (.A1(_02765_),
    .A2(\u_arbiter.i_wb_cpu_rdt[25] ),
    .ZN(_03950_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08376_ (.A1(_01437_),
    .A2(\u_arbiter.i_wb_cpu_rdt[9] ),
    .ZN(_03951_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08377_ (.A1(_03816_),
    .A2(_03950_),
    .A3(_03951_),
    .ZN(_03952_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08378_ (.A1(\u_cpu.cpu.immdec.imm30_25[1] ),
    .A2(_03740_),
    .B(_03949_),
    .C(_03952_),
    .ZN(_03953_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08379_ (.A1(_03797_),
    .A2(_03948_),
    .Z(_03954_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08380_ (.A1(\u_cpu.cpu.immdec.imm30_25[0] ),
    .A2(_03954_),
    .ZN(_03955_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08381_ (.A1(_03946_),
    .A2(_03953_),
    .B(_03955_),
    .ZN(_00909_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08382_ (.A1(_02768_),
    .A2(_03948_),
    .ZN(_03956_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08383_ (.A1(\u_cpu.cpu.immdec.imm30_25[1] ),
    .A2(_03954_),
    .B1(_03956_),
    .B2(\u_cpu.cpu.immdec.imm30_25[2] ),
    .ZN(_03957_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08384_ (.A1(_03913_),
    .A2(_03957_),
    .ZN(_00910_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08385_ (.A1(_03858_),
    .A2(_03943_),
    .ZN(_03958_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08386_ (.A1(_03761_),
    .A2(_03860_),
    .A3(_03941_),
    .ZN(_03959_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08387_ (.A1(_03773_),
    .A2(_03959_),
    .ZN(_03960_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08388_ (.A1(_03756_),
    .A2(_03810_),
    .B(_03958_),
    .C(_03960_),
    .ZN(_03961_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _08389_ (.A1(_03761_),
    .A2(_03860_),
    .B1(_03828_),
    .B2(_03788_),
    .C(_03800_),
    .ZN(_03962_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08390_ (.I0(\u_arbiter.i_wb_cpu_rdt[27] ),
    .I1(\u_arbiter.i_wb_cpu_rdt[11] ),
    .S(_01437_),
    .Z(_03963_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _08391_ (.A1(_03788_),
    .A2(_03896_),
    .B1(_03963_),
    .B2(_03779_),
    .C(_03851_),
    .ZN(_03964_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _08392_ (.A1(_03812_),
    .A2(_03961_),
    .A3(_03962_),
    .A4(_03964_),
    .Z(_03965_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _08393_ (.A1(\u_cpu.cpu.immdec.imm30_25[2] ),
    .A2(_03954_),
    .B1(_03956_),
    .B2(\u_cpu.cpu.immdec.imm30_25[3] ),
    .C1(_03963_),
    .C2(_03816_),
    .ZN(_03966_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08394_ (.A1(_03965_),
    .A2(_03966_),
    .ZN(_00911_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08395_ (.A1(_01437_),
    .A2(\u_arbiter.i_wb_cpu_rdt[12] ),
    .Z(_03967_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08396_ (.A1(_02765_),
    .A2(\u_arbiter.i_wb_cpu_rdt[28] ),
    .B(_03967_),
    .ZN(_03968_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08397_ (.A1(_03762_),
    .A2(_03891_),
    .B(_03894_),
    .ZN(_03969_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _08398_ (.A1(_03743_),
    .A2(_03786_),
    .B1(_03828_),
    .B2(_03831_),
    .C(_03904_),
    .ZN(_03970_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08399_ (.A1(_03969_),
    .A2(_03970_),
    .B(_03906_),
    .ZN(_03971_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08400_ (.A1(_01436_),
    .A2(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[9] ),
    .Z(_03972_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08401_ (.A1(_02765_),
    .A2(\u_arbiter.i_wb_cpu_rdt[9] ),
    .B(_03972_),
    .ZN(_03973_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _08402_ (.A1(_03973_),
    .A2(_03851_),
    .A3(_03826_),
    .ZN(_03974_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _08403_ (.A1(_03812_),
    .A2(_03971_),
    .A3(_03974_),
    .ZN(_03975_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08404_ (.A1(_02305_),
    .A2(_03796_),
    .A3(_03947_),
    .ZN(_03976_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _08405_ (.A1(\u_cpu.cpu.immdec.imm30_25[3] ),
    .A2(_03949_),
    .B1(_03976_),
    .B2(\u_cpu.cpu.immdec.imm30_25[4] ),
    .ZN(_03977_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08406_ (.A1(_03816_),
    .A2(_03968_),
    .B(_03975_),
    .C(_03977_),
    .ZN(_00912_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08407_ (.A1(_01437_),
    .A2(\u_arbiter.i_wb_cpu_rdt[13] ),
    .Z(_03978_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08408_ (.A1(_02765_),
    .A2(\u_arbiter.i_wb_cpu_rdt[29] ),
    .B(_03978_),
    .ZN(_03979_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08409_ (.A1(_03776_),
    .A2(_03851_),
    .ZN(_03980_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08410_ (.A1(_03742_),
    .A2(_03786_),
    .B(_03902_),
    .C(_03899_),
    .ZN(_03981_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08411_ (.A1(_03897_),
    .A2(_03981_),
    .B(_03906_),
    .ZN(_03982_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08412_ (.A1(_03927_),
    .A2(_03980_),
    .B(_03982_),
    .C(_03853_),
    .ZN(_03983_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _08413_ (.A1(\u_cpu.cpu.immdec.imm30_25[4] ),
    .A2(_03949_),
    .B1(_03976_),
    .B2(\u_cpu.cpu.immdec.imm30_25[5] ),
    .ZN(_03984_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08414_ (.A1(_03816_),
    .A2(_03979_),
    .B(_03983_),
    .C(_03984_),
    .ZN(_00913_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08415_ (.I0(\u_arbiter.i_wb_cpu_rdt[30] ),
    .I1(\u_arbiter.i_wb_cpu_rdt[14] ),
    .S(_01437_),
    .Z(_03985_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08416_ (.A1(_03742_),
    .A2(_03751_),
    .B(_03741_),
    .ZN(_03986_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _08417_ (.A1(_03741_),
    .A2(_03742_),
    .B1(_03841_),
    .B2(_03986_),
    .C(_03818_),
    .ZN(_03987_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08418_ (.A1(_03802_),
    .A2(_03826_),
    .ZN(_03988_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08419_ (.A1(_03788_),
    .A2(_03786_),
    .B(_03988_),
    .C(_03899_),
    .ZN(_03989_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08420_ (.A1(_03987_),
    .A2(_03989_),
    .B(_03906_),
    .ZN(_03990_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08421_ (.A1(_03816_),
    .A2(_03985_),
    .B1(_03990_),
    .B2(_02768_),
    .ZN(_03991_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08422_ (.A1(\u_cpu.cpu.immdec.imm30_25[5] ),
    .A2(_03954_),
    .ZN(_03992_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08423_ (.I(\u_cpu.cpu.immdec.imm19_12_20[0] ),
    .ZN(_03993_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08424_ (.A1(_01372_),
    .A2(_02313_),
    .B(\u_cpu.cpu.decode.opcode[1] ),
    .ZN(_03994_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08425_ (.A1(_02392_),
    .A2(_03994_),
    .ZN(_03995_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08426_ (.A1(_03993_),
    .A2(_03994_),
    .B(_03995_),
    .C(_02438_),
    .ZN(_03996_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08427_ (.A1(\u_cpu.cpu.immdec.imm7 ),
    .A2(_02438_),
    .B(_03956_),
    .C(_03996_),
    .ZN(_03997_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08428_ (.A1(_03991_),
    .A2(_03992_),
    .A3(_03997_),
    .ZN(_00914_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08429_ (.A1(_01436_),
    .A2(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[7] ),
    .Z(_03998_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08430_ (.A1(_02765_),
    .A2(\u_arbiter.i_wb_cpu_rdt[7] ),
    .B(_03998_),
    .ZN(_03999_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08431_ (.A1(_03807_),
    .A2(_03809_),
    .ZN(_04000_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08432_ (.A1(_03749_),
    .A2(_03831_),
    .A3(_03770_),
    .ZN(_04001_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08433_ (.A1(_03999_),
    .A2(_04000_),
    .B(_04001_),
    .C(_03755_),
    .ZN(_04002_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08434_ (.A1(_03831_),
    .A2(_03828_),
    .ZN(_04003_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08435_ (.A1(_03999_),
    .A2(_03776_),
    .ZN(_04004_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08436_ (.A1(_03744_),
    .A2(_03818_),
    .B1(_04004_),
    .B2(_03778_),
    .ZN(_04005_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _08437_ (.A1(_03999_),
    .A2(_03988_),
    .B1(_04003_),
    .B2(_04005_),
    .C(_03801_),
    .ZN(_04006_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08438_ (.A1(_03754_),
    .A2(_04002_),
    .B(_04006_),
    .ZN(_04007_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _08439_ (.A1(_03763_),
    .A2(_03778_),
    .B1(_03779_),
    .B2(_03744_),
    .C(_03851_),
    .ZN(_04008_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08440_ (.A1(_04007_),
    .A2(_04008_),
    .ZN(_04009_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08441_ (.A1(_03744_),
    .A2(_03816_),
    .B1(_04009_),
    .B2(_03876_),
    .ZN(_04010_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08442_ (.A1(_02433_),
    .A2(_02392_),
    .B(_03797_),
    .ZN(_04011_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08443_ (.A1(\u_cpu.cpu.immdec.imm7 ),
    .A2(_02305_),
    .ZN(_04012_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08444_ (.A1(_04010_),
    .A2(_04011_),
    .B1(_04012_),
    .B2(_03798_),
    .ZN(_00915_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08445_ (.A1(_01373_),
    .A2(\u_cpu.cpu.decode.opcode[1] ),
    .ZN(_04013_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08446_ (.A1(_02317_),
    .A2(_02391_),
    .A3(_04013_),
    .ZN(_04014_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08447_ (.A1(_02305_),
    .A2(_04014_),
    .B(_02767_),
    .ZN(_04015_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08448_ (.I(_04015_),
    .Z(_04016_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08449_ (.A1(\u_cpu.cpu.immdec.imm19_12_20[1] ),
    .A2(_03798_),
    .B(_04016_),
    .ZN(_04017_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08450_ (.A1(_03993_),
    .A2(_04016_),
    .B1(_04017_),
    .B2(_03855_),
    .ZN(_00916_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08451_ (.I(\u_cpu.cpu.immdec.imm19_12_20[1] ),
    .ZN(_04018_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08452_ (.A1(\u_cpu.cpu.immdec.imm19_12_20[2] ),
    .A2(_03797_),
    .B(_04016_),
    .ZN(_04019_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08453_ (.A1(_04018_),
    .A2(_04016_),
    .B1(_04019_),
    .B2(_03834_),
    .ZN(_00917_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08454_ (.I(\u_cpu.cpu.immdec.imm19_12_20[2] ),
    .ZN(_04020_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08455_ (.A1(\u_cpu.cpu.immdec.imm19_12_20[3] ),
    .A2(_03797_),
    .B(_04015_),
    .ZN(_04021_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08456_ (.A1(_04020_),
    .A2(_04016_),
    .B1(_04021_),
    .B2(_03840_),
    .ZN(_00918_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08457_ (.A1(\u_cpu.cpu.immdec.imm19_12_20[3] ),
    .A2(_04016_),
    .ZN(_04022_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _08458_ (.A1(\u_cpu.cpu.csr_imm ),
    .A2(_02305_),
    .A3(_03798_),
    .A4(_04014_),
    .ZN(_04023_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08459_ (.A1(_03845_),
    .A2(_04022_),
    .A3(_04023_),
    .ZN(_00919_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08460_ (.A1(_03973_),
    .A2(_03988_),
    .B(_03801_),
    .ZN(_04024_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08461_ (.A1(_03778_),
    .A2(_03786_),
    .ZN(_04025_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _08462_ (.A1(_03751_),
    .A2(_03765_),
    .A3(_03768_),
    .Z(_04026_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _08463_ (.A1(_03825_),
    .A2(_03776_),
    .A3(_04026_),
    .ZN(_04027_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08464_ (.A1(_04024_),
    .A2(_04025_),
    .B(_04027_),
    .ZN(_04028_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08465_ (.A1(_03851_),
    .A2(_03896_),
    .ZN(_04029_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08466_ (.A1(_03835_),
    .A2(_03988_),
    .ZN(_04030_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08467_ (.A1(_03890_),
    .A2(_03790_),
    .ZN(_04031_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _08468_ (.A1(_03999_),
    .A2(_03988_),
    .B1(_04030_),
    .B2(_04031_),
    .C(_03801_),
    .ZN(_04032_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08469_ (.A1(_04029_),
    .A2(_04004_),
    .B(_04032_),
    .C(_03782_),
    .ZN(_04033_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08470_ (.A1(_03999_),
    .A2(_04028_),
    .B(_04033_),
    .ZN(_04034_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08471_ (.A1(_03768_),
    .A2(_03774_),
    .B(_04034_),
    .C(_03740_),
    .ZN(_04035_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08472_ (.A1(\u_cpu.cpu.immdec.imm19_12_20[5] ),
    .A2(_03798_),
    .B(_04016_),
    .ZN(_04036_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08473_ (.A1(_01390_),
    .A2(_04016_),
    .B1(_04035_),
    .B2(_04036_),
    .ZN(_00920_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08474_ (.I0(\u_arbiter.i_wb_cpu_rdt[16] ),
    .I1(\u_arbiter.i_wb_cpu_rdt[0] ),
    .S(_01436_),
    .Z(_04037_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08475_ (.A1(_03779_),
    .A2(_04037_),
    .ZN(_04038_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08476_ (.A1(_03788_),
    .A2(_03776_),
    .B(_03851_),
    .C(_03896_),
    .ZN(_04039_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08477_ (.A1(_03747_),
    .A2(_03988_),
    .B(_03801_),
    .ZN(_04040_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08478_ (.A1(_03756_),
    .A2(_03789_),
    .B(_03892_),
    .ZN(_04041_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08479_ (.A1(_03828_),
    .A2(_03818_),
    .B(_03788_),
    .ZN(_04042_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08480_ (.A1(_04030_),
    .A2(_04041_),
    .A3(_04042_),
    .ZN(_04043_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _08481_ (.A1(_03747_),
    .A2(_03825_),
    .A3(_04026_),
    .B(_03851_),
    .ZN(_04044_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08482_ (.A1(_04040_),
    .A2(_04043_),
    .B(_04044_),
    .C(_03940_),
    .ZN(_04045_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08483_ (.A1(_04038_),
    .A2(_04039_),
    .B(_03782_),
    .C(_04045_),
    .ZN(_04046_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08484_ (.A1(_03782_),
    .A2(_04037_),
    .B(_04046_),
    .C(_03797_),
    .ZN(_04047_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08485_ (.A1(\u_cpu.cpu.immdec.imm19_12_20[6] ),
    .A2(_02768_),
    .ZN(_04048_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08486_ (.A1(\u_cpu.cpu.immdec.imm19_12_20[5] ),
    .A2(_04016_),
    .ZN(_04049_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _08487_ (.A1(_04016_),
    .A2(_04047_),
    .A3(_04048_),
    .B(_04049_),
    .ZN(_00921_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08488_ (.I0(\u_arbiter.i_wb_cpu_rdt[17] ),
    .I1(\u_arbiter.i_wb_cpu_rdt[1] ),
    .S(_01436_),
    .Z(_04050_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _08489_ (.A1(_03743_),
    .A2(_03776_),
    .B1(_03779_),
    .B2(_04050_),
    .C(_03851_),
    .ZN(_04051_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08490_ (.A1(_03782_),
    .A2(_04051_),
    .ZN(_04052_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08491_ (.A1(_03849_),
    .A2(_03897_),
    .ZN(_04053_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08492_ (.A1(_04024_),
    .A2(_04053_),
    .ZN(_04054_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08493_ (.A1(_03973_),
    .A2(_04028_),
    .B(_04054_),
    .C(_03851_),
    .ZN(_04055_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _08494_ (.A1(_03782_),
    .A2(_04050_),
    .B1(_04052_),
    .B2(_04055_),
    .C(_03797_),
    .ZN(_04056_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08495_ (.A1(\u_cpu.cpu.immdec.imm19_12_20[7] ),
    .A2(_02768_),
    .ZN(_04057_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08496_ (.A1(\u_cpu.cpu.immdec.imm19_12_20[6] ),
    .A2(_04016_),
    .ZN(_04058_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _08497_ (.A1(_04016_),
    .A2(_04056_),
    .A3(_04057_),
    .B(_04058_),
    .ZN(_00922_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08498_ (.I0(\u_arbiter.i_wb_cpu_rdt[18] ),
    .I1(\u_arbiter.i_wb_cpu_rdt[2] ),
    .S(_01437_),
    .Z(_04059_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08499_ (.A1(_03742_),
    .A2(_04027_),
    .B(_03780_),
    .ZN(_04060_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08500_ (.A1(_03786_),
    .A2(_03860_),
    .B(_03849_),
    .ZN(_04061_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08501_ (.A1(_03742_),
    .A2(_03897_),
    .B(_04061_),
    .C(_03791_),
    .ZN(_04062_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08502_ (.A1(_04060_),
    .A2(_04062_),
    .B(_03980_),
    .ZN(_04063_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08503_ (.A1(_03782_),
    .A2(_04059_),
    .B(_04063_),
    .C(_03797_),
    .ZN(_04064_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08504_ (.A1(\u_cpu.cpu.immdec.imm19_12_20[8] ),
    .A2(_02768_),
    .ZN(_04065_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08505_ (.A1(\u_cpu.cpu.immdec.imm19_12_20[7] ),
    .A2(_04016_),
    .ZN(_04066_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _08506_ (.A1(_04016_),
    .A2(_04064_),
    .A3(_04065_),
    .B(_04066_),
    .ZN(_00923_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08507_ (.A1(_03741_),
    .A2(_03988_),
    .ZN(_04067_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08508_ (.A1(_03849_),
    .A2(_04067_),
    .ZN(_04068_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08509_ (.A1(_01437_),
    .A2(_03668_),
    .ZN(_04069_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08510_ (.A1(_01437_),
    .A2(\u_arbiter.i_wb_cpu_rdt[19] ),
    .B(_03782_),
    .C(_04069_),
    .ZN(_04070_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08511_ (.A1(_02768_),
    .A2(_04070_),
    .ZN(_04071_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _08512_ (.A1(_03741_),
    .A2(_04027_),
    .B1(_04068_),
    .B2(_03791_),
    .C(_04071_),
    .ZN(_04072_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08513_ (.A1(_01375_),
    .A2(\u_cpu.cpu.immdec.imm24_20[0] ),
    .ZN(_04073_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08514_ (.A1(_03797_),
    .A2(_04073_),
    .ZN(_04074_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08515_ (.A1(_01374_),
    .A2(_02392_),
    .B(_04074_),
    .ZN(_04075_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08516_ (.A1(\u_cpu.cpu.immdec.imm19_12_20[8] ),
    .A2(_04016_),
    .ZN(_04076_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _08517_ (.A1(_04016_),
    .A2(_04072_),
    .A3(_04075_),
    .B(_04076_),
    .ZN(_00924_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _08518_ (.A1(_03835_),
    .A2(_03988_),
    .A3(_03902_),
    .A4(_03899_),
    .ZN(_04077_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08519_ (.I0(\u_arbiter.i_wb_cpu_rdt[31] ),
    .I1(\u_arbiter.i_wb_cpu_rdt[15] ),
    .S(_01437_),
    .Z(_04078_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08520_ (.A1(\u_cpu.cpu.immdec.imm31 ),
    .A2(_03798_),
    .B1(_03816_),
    .B2(_04078_),
    .ZN(_04079_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _08521_ (.A1(_03798_),
    .A2(_03906_),
    .A3(_04077_),
    .B(_04079_),
    .ZN(_00925_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08522_ (.I(\u_cpu.cpu.genblk3.csr.timer_irq_r ),
    .ZN(_04080_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08523_ (.A1(_02311_),
    .A2(_02448_),
    .Z(_04081_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _08524_ (.A1(\u_cpu.cpu.genblk3.csr.mie_mtie ),
    .A2(\u_cpu.cpu.genblk3.csr.mstatus_mie ),
    .A3(\u_cpu.cpu.genblk3.csr.i_mtip ),
    .A4(_04081_),
    .ZN(_04082_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08525_ (.A1(_04080_),
    .A2(_04081_),
    .B(_04082_),
    .ZN(_00926_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08526_ (.A1(_02612_),
    .A2(_02639_),
    .ZN(_04083_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08527_ (.I(_04083_),
    .Z(_04084_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08528_ (.A1(\u_cpu.rf_ram.memory[32][0] ),
    .A2(_04084_),
    .ZN(_04085_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08529_ (.A1(_03539_),
    .A2(_04084_),
    .B(_04085_),
    .ZN(_00927_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08530_ (.A1(\u_cpu.rf_ram.memory[32][1] ),
    .A2(_04084_),
    .ZN(_04086_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08531_ (.A1(_03543_),
    .A2(_04084_),
    .B(_04086_),
    .ZN(_00928_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08532_ (.A1(\u_cpu.rf_ram.memory[32][2] ),
    .A2(_04084_),
    .ZN(_04087_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08533_ (.A1(_03545_),
    .A2(_04084_),
    .B(_04087_),
    .ZN(_00929_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08534_ (.A1(\u_cpu.rf_ram.memory[32][3] ),
    .A2(_04084_),
    .ZN(_04088_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08535_ (.A1(_03547_),
    .A2(_04084_),
    .B(_04088_),
    .ZN(_00930_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08536_ (.A1(\u_cpu.rf_ram.memory[32][4] ),
    .A2(_04084_),
    .ZN(_04089_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08537_ (.A1(_03549_),
    .A2(_04084_),
    .B(_04089_),
    .ZN(_00931_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08538_ (.A1(\u_cpu.rf_ram.memory[32][5] ),
    .A2(_04084_),
    .ZN(_04090_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08539_ (.A1(_03551_),
    .A2(_04084_),
    .B(_04090_),
    .ZN(_00932_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08540_ (.A1(\u_cpu.rf_ram.memory[32][6] ),
    .A2(_04084_),
    .ZN(_04091_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08541_ (.A1(_03553_),
    .A2(_04084_),
    .B(_04091_),
    .ZN(_00933_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08542_ (.A1(\u_cpu.rf_ram.memory[32][7] ),
    .A2(_04084_),
    .ZN(_04092_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08543_ (.A1(_03555_),
    .A2(_04084_),
    .B(_04092_),
    .ZN(_00934_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08544_ (.A1(_02528_),
    .A2(_02727_),
    .ZN(_04093_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08545_ (.I(_04093_),
    .Z(_04094_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08546_ (.A1(\u_cpu.rf_ram.memory[31][0] ),
    .A2(_04094_),
    .ZN(_04095_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08547_ (.A1(_03539_),
    .A2(_04094_),
    .B(_04095_),
    .ZN(_00935_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08548_ (.A1(\u_cpu.rf_ram.memory[31][1] ),
    .A2(_04094_),
    .ZN(_04096_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08549_ (.A1(_03543_),
    .A2(_04094_),
    .B(_04096_),
    .ZN(_00936_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08550_ (.A1(\u_cpu.rf_ram.memory[31][2] ),
    .A2(_04094_),
    .ZN(_04097_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08551_ (.A1(_03545_),
    .A2(_04094_),
    .B(_04097_),
    .ZN(_00937_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08552_ (.A1(\u_cpu.rf_ram.memory[31][3] ),
    .A2(_04094_),
    .ZN(_04098_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08553_ (.A1(_03547_),
    .A2(_04094_),
    .B(_04098_),
    .ZN(_00938_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08554_ (.A1(\u_cpu.rf_ram.memory[31][4] ),
    .A2(_04094_),
    .ZN(_04099_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08555_ (.A1(_03549_),
    .A2(_04094_),
    .B(_04099_),
    .ZN(_00939_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08556_ (.A1(\u_cpu.rf_ram.memory[31][5] ),
    .A2(_04094_),
    .ZN(_04100_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08557_ (.A1(_03551_),
    .A2(_04094_),
    .B(_04100_),
    .ZN(_00940_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08558_ (.A1(\u_cpu.rf_ram.memory[31][6] ),
    .A2(_04094_),
    .ZN(_04101_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08559_ (.A1(_03553_),
    .A2(_04094_),
    .B(_04101_),
    .ZN(_00941_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08560_ (.A1(\u_cpu.rf_ram.memory[31][7] ),
    .A2(_04094_),
    .ZN(_04102_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08561_ (.A1(_03555_),
    .A2(_04094_),
    .B(_04102_),
    .ZN(_00942_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08562_ (.A1(\u_cpu.cpu.alu.cmp_r ),
    .A2(_02433_),
    .ZN(_04103_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08563_ (.A1(_02433_),
    .A2(_03494_),
    .B(_04103_),
    .ZN(_00943_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08564_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[3] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[2] ),
    .S(_02445_),
    .Z(_04104_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08565_ (.I(_04104_),
    .Z(_00944_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08566_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[4] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[3] ),
    .S(_02445_),
    .Z(_04105_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08567_ (.I(_04105_),
    .Z(_00945_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08568_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[5] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[4] ),
    .S(_02445_),
    .Z(_04106_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08569_ (.I(_04106_),
    .Z(_00946_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08570_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[6] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[5] ),
    .S(_02445_),
    .Z(_04107_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08571_ (.I(_04107_),
    .Z(_00947_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08572_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[7] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[6] ),
    .S(_02445_),
    .Z(_04108_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08573_ (.I(_04108_),
    .Z(_00948_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08574_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[8] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[7] ),
    .S(_02445_),
    .Z(_04109_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08575_ (.I(_04109_),
    .Z(_00949_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08576_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[9] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[8] ),
    .S(_02445_),
    .Z(_04110_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08577_ (.I(_04110_),
    .Z(_00950_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08578_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[10] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[9] ),
    .S(_02445_),
    .Z(_04111_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08579_ (.I(_04111_),
    .Z(_00951_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08580_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[11] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[10] ),
    .S(_02445_),
    .Z(_04112_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08581_ (.I(_04112_),
    .Z(_00952_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08582_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[12] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[11] ),
    .S(_02445_),
    .Z(_04113_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08583_ (.I(_04113_),
    .Z(_00953_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08584_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[13] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[12] ),
    .S(_02445_),
    .Z(_04114_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08585_ (.I(_04114_),
    .Z(_00954_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08586_ (.I(_02372_),
    .Z(_04115_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08587_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[14] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[13] ),
    .S(_04115_),
    .Z(_04116_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08588_ (.I(_04116_),
    .Z(_00955_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08589_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[15] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[14] ),
    .S(_04115_),
    .Z(_04117_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08590_ (.I(_04117_),
    .Z(_00956_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08591_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[16] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[15] ),
    .S(_04115_),
    .Z(_04118_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08592_ (.I(_04118_),
    .Z(_00957_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08593_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[17] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[16] ),
    .S(_04115_),
    .Z(_04119_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08594_ (.I(_04119_),
    .Z(_00958_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08595_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[18] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[17] ),
    .S(_04115_),
    .Z(_04120_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08596_ (.I(_04120_),
    .Z(_00959_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08597_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[19] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[18] ),
    .S(_04115_),
    .Z(_04121_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08598_ (.I(_04121_),
    .Z(_00960_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08599_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[20] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[19] ),
    .S(_04115_),
    .Z(_04122_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08600_ (.I(_04122_),
    .Z(_00961_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08601_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[21] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[20] ),
    .S(_04115_),
    .Z(_04123_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08602_ (.I(_04123_),
    .Z(_00962_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08603_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[22] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[21] ),
    .S(_04115_),
    .Z(_04124_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08604_ (.I(_04124_),
    .Z(_00963_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08605_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[23] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[22] ),
    .S(_04115_),
    .Z(_04125_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08606_ (.I(_04125_),
    .Z(_00964_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08607_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[24] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[23] ),
    .S(_04115_),
    .Z(_04126_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08608_ (.I(_04126_),
    .Z(_00965_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08609_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[25] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[24] ),
    .S(_04115_),
    .Z(_04127_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08610_ (.I(_04127_),
    .Z(_00966_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08611_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[26] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[25] ),
    .S(_04115_),
    .Z(_04128_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08612_ (.I(_04128_),
    .Z(_00967_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08613_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[27] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[26] ),
    .S(_04115_),
    .Z(_04129_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08614_ (.I(_04129_),
    .Z(_00968_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08615_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[28] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[27] ),
    .S(_04115_),
    .Z(_04130_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08616_ (.I(_04130_),
    .Z(_00969_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08617_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[29] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[28] ),
    .S(_04115_),
    .Z(_04131_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08618_ (.I(_04131_),
    .Z(_00970_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08619_ (.I0(\u_arbiter.i_wb_cpu_dbus_adr[30] ),
    .I1(\u_arbiter.i_wb_cpu_dbus_adr[29] ),
    .S(_02372_),
    .Z(_04132_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08620_ (.I(_04132_),
    .Z(_00971_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08621_ (.I(\u_arbiter.i_wb_cpu_dbus_adr[31] ),
    .ZN(_04133_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08622_ (.A1(\u_arbiter.i_wb_cpu_dbus_adr[30] ),
    .A2(_02445_),
    .ZN(_04134_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08623_ (.A1(_04133_),
    .A2(_02445_),
    .B(_04134_),
    .ZN(_00972_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08624_ (.A1(\u_cpu.cpu.bufreg.i_sh_signed ),
    .A2(_02448_),
    .B(_02445_),
    .ZN(_04135_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _08625_ (.A1(_01372_),
    .A2(_02394_),
    .A3(_02441_),
    .B(_02443_),
    .ZN(_04136_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08626_ (.A1(_02444_),
    .A2(_02773_),
    .A3(_04136_),
    .ZN(_04137_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _08627_ (.A1(_04133_),
    .A2(_04135_),
    .B1(_04137_),
    .B2(_02445_),
    .ZN(_00973_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08628_ (.A1(\u_cpu.cpu.state.o_cnt_r[0] ),
    .A2(\u_cpu.cpu.state.o_cnt_r[1] ),
    .B(_02338_),
    .C(_02773_),
    .ZN(_04138_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08629_ (.A1(_02372_),
    .A2(_02773_),
    .B(_04138_),
    .ZN(_04139_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08630_ (.A1(\u_cpu.cpu.bufreg.lsb[1] ),
    .A2(_04139_),
    .ZN(_04140_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08631_ (.A1(_02361_),
    .A2(_04139_),
    .B(_04140_),
    .ZN(_00974_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08632_ (.A1(\u_arbiter.i_wb_cpu_dbus_adr[2] ),
    .A2(_02448_),
    .ZN(_04141_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08633_ (.A1(_04137_),
    .A2(_04141_),
    .ZN(_04142_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08634_ (.A1(_04139_),
    .A2(_04142_),
    .ZN(_04143_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08635_ (.A1(_02431_),
    .A2(_04139_),
    .B(_04143_),
    .ZN(_00975_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08636_ (.A1(_02528_),
    .A2(_02625_),
    .ZN(_04144_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08637_ (.I(_04144_),
    .Z(_04145_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08638_ (.A1(\u_cpu.rf_ram.memory[30][0] ),
    .A2(_04145_),
    .ZN(_04146_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08639_ (.A1(_03539_),
    .A2(_04145_),
    .B(_04146_),
    .ZN(_00976_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08640_ (.A1(\u_cpu.rf_ram.memory[30][1] ),
    .A2(_04145_),
    .ZN(_04147_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08641_ (.A1(_03543_),
    .A2(_04145_),
    .B(_04147_),
    .ZN(_00977_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08642_ (.A1(\u_cpu.rf_ram.memory[30][2] ),
    .A2(_04145_),
    .ZN(_04148_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08643_ (.A1(_03545_),
    .A2(_04145_),
    .B(_04148_),
    .ZN(_00978_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08644_ (.A1(\u_cpu.rf_ram.memory[30][3] ),
    .A2(_04145_),
    .ZN(_04149_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08645_ (.A1(_03547_),
    .A2(_04145_),
    .B(_04149_),
    .ZN(_00979_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08646_ (.A1(\u_cpu.rf_ram.memory[30][4] ),
    .A2(_04145_),
    .ZN(_04150_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08647_ (.A1(_03549_),
    .A2(_04145_),
    .B(_04150_),
    .ZN(_00980_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08648_ (.A1(\u_cpu.rf_ram.memory[30][5] ),
    .A2(_04145_),
    .ZN(_04151_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08649_ (.A1(_03551_),
    .A2(_04145_),
    .B(_04151_),
    .ZN(_00981_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08650_ (.A1(\u_cpu.rf_ram.memory[30][6] ),
    .A2(_04145_),
    .ZN(_04152_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08651_ (.A1(_03553_),
    .A2(_04145_),
    .B(_04152_),
    .ZN(_00982_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08652_ (.A1(\u_cpu.rf_ram.memory[30][7] ),
    .A2(_04145_),
    .ZN(_04153_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08653_ (.A1(_03555_),
    .A2(_04145_),
    .B(_04153_),
    .ZN(_00983_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08654_ (.A1(_02305_),
    .A2(_02448_),
    .B(_01428_),
    .ZN(_04154_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08655_ (.I(_04154_),
    .Z(_04155_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08656_ (.A1(_01428_),
    .A2(_02449_),
    .ZN(_04156_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08657_ (.I(_04156_),
    .Z(_04157_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08658_ (.A1(\u_arbiter.i_wb_cpu_ibus_adr[0] ),
    .A2(_04155_),
    .B1(_04157_),
    .B2(\u_arbiter.i_wb_cpu_ibus_adr[1] ),
    .ZN(_04158_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _08659_ (.I(_04158_),
    .ZN(_00984_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08660_ (.A1(\u_arbiter.i_wb_cpu_ibus_adr[1] ),
    .A2(_04155_),
    .B1(_04157_),
    .B2(\u_cpu.cpu.ctrl.o_ibus_adr[2] ),
    .ZN(_04159_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _08661_ (.I(_04159_),
    .ZN(_00985_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08662_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[2] ),
    .A2(_04155_),
    .B1(_04157_),
    .B2(\u_cpu.cpu.ctrl.o_ibus_adr[3] ),
    .ZN(_04160_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _08663_ (.I(_04160_),
    .ZN(_00986_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08664_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[3] ),
    .A2(_04155_),
    .B1(_04157_),
    .B2(\u_cpu.cpu.ctrl.o_ibus_adr[4] ),
    .ZN(_04161_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _08665_ (.I(_04161_),
    .ZN(_00987_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08666_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[4] ),
    .A2(_04155_),
    .B1(_04157_),
    .B2(\u_cpu.cpu.ctrl.o_ibus_adr[5] ),
    .ZN(_04162_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _08667_ (.I(_04162_),
    .ZN(_00988_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08668_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[5] ),
    .A2(_04155_),
    .B1(_04157_),
    .B2(\u_cpu.cpu.ctrl.o_ibus_adr[6] ),
    .ZN(_04163_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _08669_ (.I(_04163_),
    .ZN(_00989_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08670_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[6] ),
    .A2(_04155_),
    .B1(_04157_),
    .B2(\u_cpu.cpu.ctrl.o_ibus_adr[7] ),
    .ZN(_04164_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _08671_ (.I(_04164_),
    .ZN(_00990_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08672_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[7] ),
    .A2(_04155_),
    .B1(_04157_),
    .B2(\u_cpu.cpu.ctrl.o_ibus_adr[8] ),
    .ZN(_04165_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _08673_ (.I(_04165_),
    .ZN(_00991_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08674_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[8] ),
    .A2(_04155_),
    .B1(_04157_),
    .B2(\u_cpu.cpu.ctrl.o_ibus_adr[9] ),
    .ZN(_04166_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _08675_ (.I(_04166_),
    .ZN(_00992_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08676_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[9] ),
    .A2(_04155_),
    .B1(_04157_),
    .B2(\u_cpu.cpu.ctrl.o_ibus_adr[10] ),
    .ZN(_04167_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _08677_ (.I(_04167_),
    .ZN(_00993_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08678_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[10] ),
    .A2(_04155_),
    .B1(_04157_),
    .B2(\u_cpu.cpu.ctrl.o_ibus_adr[11] ),
    .ZN(_04168_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _08679_ (.I(_04168_),
    .ZN(_00994_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08680_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[11] ),
    .A2(_04155_),
    .B1(_04157_),
    .B2(\u_cpu.cpu.ctrl.o_ibus_adr[12] ),
    .ZN(_04169_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _08681_ (.I(_04169_),
    .ZN(_00995_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08682_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[12] ),
    .A2(_04155_),
    .B1(_04157_),
    .B2(\u_cpu.cpu.ctrl.o_ibus_adr[13] ),
    .ZN(_04170_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _08683_ (.I(_04170_),
    .ZN(_00996_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08684_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[13] ),
    .A2(_04155_),
    .B1(_04157_),
    .B2(\u_cpu.cpu.ctrl.o_ibus_adr[14] ),
    .ZN(_04171_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _08685_ (.I(_04171_),
    .ZN(_00997_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08686_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[14] ),
    .A2(_04155_),
    .B1(_04157_),
    .B2(\u_cpu.cpu.ctrl.o_ibus_adr[15] ),
    .ZN(_04172_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _08687_ (.I(_04172_),
    .ZN(_00998_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08688_ (.I(_04154_),
    .Z(_04173_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08689_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[15] ),
    .A2(_04173_),
    .B1(_04157_),
    .B2(\u_cpu.cpu.ctrl.o_ibus_adr[16] ),
    .ZN(_04174_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _08690_ (.I(_04174_),
    .ZN(_00999_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08691_ (.I(_04156_),
    .Z(_04175_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08692_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[16] ),
    .A2(_04173_),
    .B1(_04175_),
    .B2(\u_cpu.cpu.ctrl.o_ibus_adr[17] ),
    .ZN(_04176_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _08693_ (.I(_04176_),
    .ZN(_01000_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08694_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[17] ),
    .A2(_04173_),
    .B1(_04175_),
    .B2(\u_cpu.cpu.ctrl.o_ibus_adr[18] ),
    .ZN(_04177_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _08695_ (.I(_04177_),
    .ZN(_01001_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08696_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[18] ),
    .A2(_04173_),
    .B1(_04175_),
    .B2(\u_cpu.cpu.ctrl.o_ibus_adr[19] ),
    .ZN(_04178_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _08697_ (.I(_04178_),
    .ZN(_01002_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08698_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[19] ),
    .A2(_04173_),
    .B1(_04175_),
    .B2(\u_cpu.cpu.ctrl.o_ibus_adr[20] ),
    .ZN(_04179_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _08699_ (.I(_04179_),
    .ZN(_01003_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08700_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[20] ),
    .A2(_04173_),
    .B1(_04175_),
    .B2(\u_cpu.cpu.ctrl.o_ibus_adr[21] ),
    .ZN(_04180_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _08701_ (.I(_04180_),
    .ZN(_01004_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08702_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[21] ),
    .A2(_04173_),
    .B1(_04175_),
    .B2(\u_cpu.cpu.ctrl.o_ibus_adr[22] ),
    .ZN(_04181_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _08703_ (.I(_04181_),
    .ZN(_01005_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08704_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[22] ),
    .A2(_04173_),
    .B1(_04175_),
    .B2(\u_cpu.cpu.ctrl.o_ibus_adr[23] ),
    .ZN(_04182_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _08705_ (.I(_04182_),
    .ZN(_01006_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08706_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[23] ),
    .A2(_04173_),
    .B1(_04175_),
    .B2(\u_cpu.cpu.ctrl.o_ibus_adr[24] ),
    .ZN(_04183_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _08707_ (.I(_04183_),
    .ZN(_01007_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08708_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[24] ),
    .A2(_04173_),
    .B1(_04175_),
    .B2(\u_cpu.cpu.ctrl.o_ibus_adr[25] ),
    .ZN(_04184_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _08709_ (.I(_04184_),
    .ZN(_01008_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08710_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[25] ),
    .A2(_04173_),
    .B1(_04175_),
    .B2(\u_cpu.cpu.ctrl.o_ibus_adr[26] ),
    .ZN(_04185_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _08711_ (.I(_04185_),
    .ZN(_01009_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08712_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[26] ),
    .A2(_04173_),
    .B1(_04175_),
    .B2(\u_cpu.cpu.ctrl.o_ibus_adr[27] ),
    .ZN(_04186_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _08713_ (.I(_04186_),
    .ZN(_01010_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08714_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[27] ),
    .A2(_04173_),
    .B1(_04175_),
    .B2(\u_cpu.cpu.ctrl.o_ibus_adr[28] ),
    .ZN(_04187_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _08715_ (.I(_04187_),
    .ZN(_01011_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08716_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[28] ),
    .A2(_04173_),
    .B1(_04175_),
    .B2(\u_cpu.cpu.ctrl.o_ibus_adr[29] ),
    .ZN(_04188_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _08717_ (.I(_04188_),
    .ZN(_01012_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08718_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[29] ),
    .A2(_04173_),
    .B1(_04175_),
    .B2(\u_cpu.cpu.ctrl.o_ibus_adr[30] ),
    .ZN(_04189_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _08719_ (.I(_04189_),
    .ZN(_01013_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08720_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[30] ),
    .A2(_04173_),
    .B1(_04175_),
    .B2(\u_cpu.cpu.ctrl.o_ibus_adr[31] ),
    .ZN(_04190_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _08721_ (.I(_04190_),
    .ZN(_01014_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _08722_ (.A1(_02343_),
    .A2(_01410_),
    .A3(_01378_),
    .ZN(_04191_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08723_ (.A1(_04191_),
    .A2(_01386_),
    .ZN(_04192_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08724_ (.I0(_02381_),
    .I1(_02406_),
    .S(\u_cpu.cpu.ctrl.i_jump ),
    .Z(_04193_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08725_ (.A1(_02324_),
    .A2(_02356_),
    .B(_04192_),
    .ZN(_04194_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08726_ (.A1(_04192_),
    .A2(_04193_),
    .B(_04194_),
    .ZN(_04195_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08727_ (.A1(\u_cpu.cpu.ctrl.o_ibus_adr[31] ),
    .A2(_04154_),
    .B1(_04175_),
    .B2(_04195_),
    .ZN(_04196_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _08728_ (.I(_04196_),
    .ZN(_01015_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _08729_ (.A1(\u_cpu.cpu.immdec.imm11_7[2] ),
    .A2(_02473_),
    .A3(_02574_),
    .ZN(_04197_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08730_ (.A1(_02660_),
    .A2(_04197_),
    .ZN(_04198_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08731_ (.I(_04198_),
    .Z(_04199_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08732_ (.A1(\u_cpu.rf_ram.memory[109][0] ),
    .A2(_04199_),
    .ZN(_04200_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08733_ (.A1(_03539_),
    .A2(_04199_),
    .B(_04200_),
    .ZN(_01016_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08734_ (.A1(\u_cpu.rf_ram.memory[109][1] ),
    .A2(_04199_),
    .ZN(_04201_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08735_ (.A1(_03543_),
    .A2(_04199_),
    .B(_04201_),
    .ZN(_01017_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08736_ (.A1(\u_cpu.rf_ram.memory[109][2] ),
    .A2(_04199_),
    .ZN(_04202_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08737_ (.A1(_03545_),
    .A2(_04199_),
    .B(_04202_),
    .ZN(_01018_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08738_ (.A1(\u_cpu.rf_ram.memory[109][3] ),
    .A2(_04199_),
    .ZN(_04203_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08739_ (.A1(_03547_),
    .A2(_04199_),
    .B(_04203_),
    .ZN(_01019_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08740_ (.A1(\u_cpu.rf_ram.memory[109][4] ),
    .A2(_04199_),
    .ZN(_04204_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08741_ (.A1(_03549_),
    .A2(_04199_),
    .B(_04204_),
    .ZN(_01020_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08742_ (.A1(\u_cpu.rf_ram.memory[109][5] ),
    .A2(_04199_),
    .ZN(_04205_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08743_ (.A1(_03551_),
    .A2(_04199_),
    .B(_04205_),
    .ZN(_01021_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08744_ (.A1(\u_cpu.rf_ram.memory[109][6] ),
    .A2(_04199_),
    .ZN(_04206_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08745_ (.A1(_03553_),
    .A2(_04199_),
    .B(_04206_),
    .ZN(_01022_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08746_ (.A1(\u_cpu.rf_ram.memory[109][7] ),
    .A2(_04199_),
    .ZN(_04207_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08747_ (.A1(_03555_),
    .A2(_04199_),
    .B(_04207_),
    .ZN(_01023_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08748_ (.A1(_02577_),
    .A2(_02682_),
    .ZN(_04208_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08749_ (.I0(_02573_),
    .I1(\u_cpu.rf_ram.memory[3][0] ),
    .S(_04208_),
    .Z(_04209_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08750_ (.I(_04209_),
    .Z(_01024_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08751_ (.I0(_02581_),
    .I1(\u_cpu.rf_ram.memory[3][1] ),
    .S(_04208_),
    .Z(_04210_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08752_ (.I(_04210_),
    .Z(_01025_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08753_ (.I0(_02584_),
    .I1(\u_cpu.rf_ram.memory[3][2] ),
    .S(_04208_),
    .Z(_04211_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08754_ (.I(_04211_),
    .Z(_01026_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08755_ (.I0(_02587_),
    .I1(\u_cpu.rf_ram.memory[3][3] ),
    .S(_04208_),
    .Z(_04212_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08756_ (.I(_04212_),
    .Z(_01027_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08757_ (.I0(_02590_),
    .I1(\u_cpu.rf_ram.memory[3][4] ),
    .S(_04208_),
    .Z(_04213_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08758_ (.I(_04213_),
    .Z(_01028_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08759_ (.I0(_02593_),
    .I1(\u_cpu.rf_ram.memory[3][5] ),
    .S(_04208_),
    .Z(_04214_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08760_ (.I(_04214_),
    .Z(_01029_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08761_ (.I0(_02596_),
    .I1(\u_cpu.rf_ram.memory[3][6] ),
    .S(_04208_),
    .Z(_04215_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08762_ (.I(_04215_),
    .Z(_01030_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08763_ (.I0(_02599_),
    .I1(\u_cpu.rf_ram.memory[3][7] ),
    .S(_04208_),
    .Z(_04216_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08764_ (.I(_04216_),
    .Z(_01031_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08765_ (.A1(_02469_),
    .A2(_02577_),
    .ZN(_04217_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08766_ (.I0(_02573_),
    .I1(\u_cpu.rf_ram.memory[2][0] ),
    .S(_04217_),
    .Z(_04218_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08767_ (.I(_04218_),
    .Z(_01032_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08768_ (.I0(_02581_),
    .I1(\u_cpu.rf_ram.memory[2][1] ),
    .S(_04217_),
    .Z(_04219_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08769_ (.I(_04219_),
    .Z(_01033_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08770_ (.I0(_02584_),
    .I1(\u_cpu.rf_ram.memory[2][2] ),
    .S(_04217_),
    .Z(_04220_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08771_ (.I(_04220_),
    .Z(_01034_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08772_ (.I0(_02587_),
    .I1(\u_cpu.rf_ram.memory[2][3] ),
    .S(_04217_),
    .Z(_04221_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08773_ (.I(_04221_),
    .Z(_01035_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08774_ (.I0(_02590_),
    .I1(\u_cpu.rf_ram.memory[2][4] ),
    .S(_04217_),
    .Z(_04222_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08775_ (.I(_04222_),
    .Z(_01036_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08776_ (.I0(_02593_),
    .I1(\u_cpu.rf_ram.memory[2][5] ),
    .S(_04217_),
    .Z(_04223_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08777_ (.I(_04223_),
    .Z(_01037_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08778_ (.I0(_02596_),
    .I1(\u_cpu.rf_ram.memory[2][6] ),
    .S(_04217_),
    .Z(_04224_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08779_ (.I(_04224_),
    .Z(_01038_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08780_ (.I0(_02599_),
    .I1(\u_cpu.rf_ram.memory[2][7] ),
    .S(_04217_),
    .Z(_04225_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08781_ (.I(_04225_),
    .Z(_01039_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08782_ (.A1(_02475_),
    .A2(_02660_),
    .ZN(_04226_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08783_ (.I(_04226_),
    .Z(_04227_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08784_ (.A1(\u_cpu.rf_ram.memory[93][0] ),
    .A2(_04227_),
    .ZN(_04228_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08785_ (.A1(_03539_),
    .A2(_04227_),
    .B(_04228_),
    .ZN(_01040_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08786_ (.A1(\u_cpu.rf_ram.memory[93][1] ),
    .A2(_04227_),
    .ZN(_04229_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08787_ (.A1(_03543_),
    .A2(_04227_),
    .B(_04229_),
    .ZN(_01041_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08788_ (.A1(\u_cpu.rf_ram.memory[93][2] ),
    .A2(_04227_),
    .ZN(_04230_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08789_ (.A1(_03545_),
    .A2(_04227_),
    .B(_04230_),
    .ZN(_01042_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08790_ (.A1(\u_cpu.rf_ram.memory[93][3] ),
    .A2(_04227_),
    .ZN(_04231_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08791_ (.A1(_03547_),
    .A2(_04227_),
    .B(_04231_),
    .ZN(_01043_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08792_ (.A1(\u_cpu.rf_ram.memory[93][4] ),
    .A2(_04227_),
    .ZN(_04232_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08793_ (.A1(_03549_),
    .A2(_04227_),
    .B(_04232_),
    .ZN(_01044_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08794_ (.A1(\u_cpu.rf_ram.memory[93][5] ),
    .A2(_04227_),
    .ZN(_04233_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08795_ (.A1(_03551_),
    .A2(_04227_),
    .B(_04233_),
    .ZN(_01045_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08796_ (.A1(\u_cpu.rf_ram.memory[93][6] ),
    .A2(_04227_),
    .ZN(_04234_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08797_ (.A1(_03553_),
    .A2(_04227_),
    .B(_04234_),
    .ZN(_01046_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08798_ (.A1(\u_cpu.rf_ram.memory[93][7] ),
    .A2(_04227_),
    .ZN(_04235_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08799_ (.A1(_03555_),
    .A2(_04227_),
    .B(_04235_),
    .ZN(_01047_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08800_ (.A1(_02433_),
    .A2(_02453_),
    .ZN(_04236_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08801_ (.A1(_02768_),
    .A2(_04236_),
    .ZN(_04237_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08802_ (.A1(\u_cpu.cpu.immdec.imm11_7[1] ),
    .A2(_03797_),
    .B(_04237_),
    .ZN(_04238_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08803_ (.A1(_02312_),
    .A2(_04237_),
    .B1(_04238_),
    .B2(_04010_),
    .ZN(_01048_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08804_ (.A1(_03860_),
    .A2(_03818_),
    .B(_03788_),
    .ZN(_04239_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08805_ (.A1(_03857_),
    .A2(_03897_),
    .A3(_04239_),
    .ZN(_04240_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08806_ (.A1(_04040_),
    .A2(_04240_),
    .B(_03780_),
    .ZN(_04241_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _08807_ (.A1(_03747_),
    .A2(_03825_),
    .A3(_04000_),
    .B1(_04241_),
    .B2(_03782_),
    .ZN(_04242_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08808_ (.A1(_03761_),
    .A2(_03778_),
    .B1(_03779_),
    .B2(_03788_),
    .ZN(_04243_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08809_ (.A1(_03780_),
    .A2(_04243_),
    .ZN(_04244_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08810_ (.A1(_03740_),
    .A2(_04242_),
    .A3(_04244_),
    .ZN(_04245_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08811_ (.I0(\u_cpu.cpu.immdec.imm11_7[1] ),
    .I1(\u_cpu.cpu.immdec.imm11_7[2] ),
    .S(_04236_),
    .Z(_04246_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08812_ (.A1(_03788_),
    .A2(_03816_),
    .B1(_04246_),
    .B2(_03798_),
    .ZN(_04247_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08813_ (.A1(_04245_),
    .A2(_04247_),
    .ZN(_01049_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08814_ (.A1(_03762_),
    .A2(_03778_),
    .ZN(_04248_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _08815_ (.A1(_03973_),
    .A2(_03769_),
    .B1(_03809_),
    .B2(_03757_),
    .C(_04248_),
    .ZN(_04249_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08816_ (.A1(_03743_),
    .A2(_03826_),
    .ZN(_04250_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08817_ (.A1(_03810_),
    .A2(_04250_),
    .B(_03897_),
    .C(_03873_),
    .ZN(_04251_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08818_ (.A1(_03780_),
    .A2(_04249_),
    .B1(_04251_),
    .B2(_04024_),
    .ZN(_04252_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08819_ (.A1(_03812_),
    .A2(_04252_),
    .ZN(_04253_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08820_ (.A1(\u_cpu.cpu.immdec.imm11_7[3] ),
    .A2(_03798_),
    .B(_04253_),
    .ZN(_04254_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08821_ (.A1(_03825_),
    .A2(_03770_),
    .ZN(_04255_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08822_ (.A1(_03782_),
    .A2(_04255_),
    .ZN(_04256_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08823_ (.A1(_03973_),
    .A2(_04256_),
    .ZN(_04257_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08824_ (.A1(\u_cpu.cpu.immdec.imm11_7[2] ),
    .A2(_04237_),
    .B1(_04257_),
    .B2(_03740_),
    .ZN(_04258_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08825_ (.A1(_04237_),
    .A2(_04254_),
    .B(_04258_),
    .ZN(_01050_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08826_ (.A1(_03755_),
    .A2(_03786_),
    .B(_04256_),
    .C(_03851_),
    .ZN(_04259_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08827_ (.A1(_03778_),
    .A2(_03780_),
    .B1(_04259_),
    .B2(_03742_),
    .ZN(_04260_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08828_ (.A1(_03801_),
    .A2(_03900_),
    .B(_04260_),
    .ZN(_04261_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08829_ (.A1(\u_cpu.cpu.immdec.imm11_7[3] ),
    .A2(_04236_),
    .ZN(_04262_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08830_ (.A1(_02525_),
    .A2(_04236_),
    .B(_04262_),
    .ZN(_04263_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08831_ (.I0(_04261_),
    .I1(_04263_),
    .S(_03797_),
    .Z(_04264_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08832_ (.I(_04264_),
    .Z(_01051_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08833_ (.A1(_03773_),
    .A2(_03787_),
    .ZN(_04265_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08834_ (.A1(_03861_),
    .A2(_04265_),
    .B(_03807_),
    .C(_03851_),
    .ZN(_04266_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08835_ (.A1(_03811_),
    .A2(_03809_),
    .A3(_04266_),
    .ZN(_04267_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08836_ (.A1(_03740_),
    .A2(_03741_),
    .A3(_04267_),
    .ZN(_04268_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08837_ (.A1(\u_cpu.cpu.immdec.imm30_25[0] ),
    .A2(_03798_),
    .B(_04237_),
    .ZN(_04269_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08838_ (.A1(_02525_),
    .A2(_04237_),
    .B1(_04268_),
    .B2(_04269_),
    .ZN(_01052_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08839_ (.A1(_02539_),
    .A2(_04197_),
    .ZN(_04270_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08840_ (.I(_04270_),
    .Z(_04271_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08841_ (.A1(\u_cpu.rf_ram.memory[97][0] ),
    .A2(_04271_),
    .ZN(_04272_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08842_ (.A1(_03539_),
    .A2(_04271_),
    .B(_04272_),
    .ZN(_01053_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08843_ (.A1(\u_cpu.rf_ram.memory[97][1] ),
    .A2(_04271_),
    .ZN(_04273_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08844_ (.A1(_03543_),
    .A2(_04271_),
    .B(_04273_),
    .ZN(_01054_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08845_ (.A1(\u_cpu.rf_ram.memory[97][2] ),
    .A2(_04271_),
    .ZN(_04274_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08846_ (.A1(_03545_),
    .A2(_04271_),
    .B(_04274_),
    .ZN(_01055_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08847_ (.A1(\u_cpu.rf_ram.memory[97][3] ),
    .A2(_04271_),
    .ZN(_04275_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08848_ (.A1(_03547_),
    .A2(_04271_),
    .B(_04275_),
    .ZN(_01056_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08849_ (.A1(\u_cpu.rf_ram.memory[97][4] ),
    .A2(_04271_),
    .ZN(_04276_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08850_ (.A1(_03549_),
    .A2(_04271_),
    .B(_04276_),
    .ZN(_01057_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08851_ (.A1(\u_cpu.rf_ram.memory[97][5] ),
    .A2(_04271_),
    .ZN(_04277_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08852_ (.A1(_03551_),
    .A2(_04271_),
    .B(_04277_),
    .ZN(_01058_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08853_ (.A1(\u_cpu.rf_ram.memory[97][6] ),
    .A2(_04271_),
    .ZN(_04278_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08854_ (.A1(_03553_),
    .A2(_04271_),
    .B(_04278_),
    .ZN(_01059_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08855_ (.A1(\u_cpu.rf_ram.memory[97][7] ),
    .A2(_04271_),
    .ZN(_04279_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08856_ (.A1(_03555_),
    .A2(_04271_),
    .B(_04279_),
    .ZN(_01060_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08857_ (.I(_02481_),
    .Z(_04280_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08858_ (.A1(_02475_),
    .A2(_02625_),
    .ZN(_04281_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08859_ (.I(_04281_),
    .Z(_04282_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08860_ (.A1(\u_cpu.rf_ram.memory[94][0] ),
    .A2(_04282_),
    .ZN(_04283_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08861_ (.A1(_04280_),
    .A2(_04282_),
    .B(_04283_),
    .ZN(_01061_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08862_ (.I(_02486_),
    .Z(_04284_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08863_ (.A1(\u_cpu.rf_ram.memory[94][1] ),
    .A2(_04282_),
    .ZN(_04285_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08864_ (.A1(_04284_),
    .A2(_04282_),
    .B(_04285_),
    .ZN(_01062_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08865_ (.I(_02491_),
    .Z(_04286_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08866_ (.A1(\u_cpu.rf_ram.memory[94][2] ),
    .A2(_04282_),
    .ZN(_04287_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08867_ (.A1(_04286_),
    .A2(_04282_),
    .B(_04287_),
    .ZN(_01063_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08868_ (.I(_02496_),
    .Z(_04288_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08869_ (.A1(\u_cpu.rf_ram.memory[94][3] ),
    .A2(_04282_),
    .ZN(_04289_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08870_ (.A1(_04288_),
    .A2(_04282_),
    .B(_04289_),
    .ZN(_01064_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08871_ (.I(_02501_),
    .Z(_04290_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08872_ (.A1(\u_cpu.rf_ram.memory[94][4] ),
    .A2(_04282_),
    .ZN(_04291_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08873_ (.A1(_04290_),
    .A2(_04282_),
    .B(_04291_),
    .ZN(_01065_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08874_ (.I(_02506_),
    .Z(_04292_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08875_ (.A1(\u_cpu.rf_ram.memory[94][5] ),
    .A2(_04282_),
    .ZN(_04293_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08876_ (.A1(_04292_),
    .A2(_04282_),
    .B(_04293_),
    .ZN(_01066_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08877_ (.I(_02511_),
    .Z(_04294_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08878_ (.A1(\u_cpu.rf_ram.memory[94][6] ),
    .A2(_04282_),
    .ZN(_04295_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08879_ (.A1(_04294_),
    .A2(_04282_),
    .B(_04295_),
    .ZN(_01067_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08880_ (.I(_02516_),
    .Z(_04296_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08881_ (.A1(\u_cpu.rf_ram.memory[94][7] ),
    .A2(_04282_),
    .ZN(_04297_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08882_ (.A1(_04296_),
    .A2(_04282_),
    .B(_04297_),
    .ZN(_01068_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08883_ (.A1(_02475_),
    .A2(_02727_),
    .ZN(_04298_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08884_ (.I(_04298_),
    .Z(_04299_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08885_ (.A1(\u_cpu.rf_ram.memory[95][0] ),
    .A2(_04299_),
    .ZN(_04300_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08886_ (.A1(_04280_),
    .A2(_04299_),
    .B(_04300_),
    .ZN(_01069_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08887_ (.A1(\u_cpu.rf_ram.memory[95][1] ),
    .A2(_04299_),
    .ZN(_04301_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08888_ (.A1(_04284_),
    .A2(_04299_),
    .B(_04301_),
    .ZN(_01070_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08889_ (.A1(\u_cpu.rf_ram.memory[95][2] ),
    .A2(_04299_),
    .ZN(_04302_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08890_ (.A1(_04286_),
    .A2(_04299_),
    .B(_04302_),
    .ZN(_01071_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08891_ (.A1(\u_cpu.rf_ram.memory[95][3] ),
    .A2(_04299_),
    .ZN(_04303_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08892_ (.A1(_04288_),
    .A2(_04299_),
    .B(_04303_),
    .ZN(_01072_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08893_ (.A1(\u_cpu.rf_ram.memory[95][4] ),
    .A2(_04299_),
    .ZN(_04304_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08894_ (.A1(_04290_),
    .A2(_04299_),
    .B(_04304_),
    .ZN(_01073_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08895_ (.A1(\u_cpu.rf_ram.memory[95][5] ),
    .A2(_04299_),
    .ZN(_04305_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08896_ (.A1(_04292_),
    .A2(_04299_),
    .B(_04305_),
    .ZN(_01074_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08897_ (.A1(\u_cpu.rf_ram.memory[95][6] ),
    .A2(_04299_),
    .ZN(_04306_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08898_ (.A1(_04294_),
    .A2(_04299_),
    .B(_04306_),
    .ZN(_01075_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08899_ (.A1(\u_cpu.rf_ram.memory[95][7] ),
    .A2(_04299_),
    .ZN(_04307_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08900_ (.A1(_04296_),
    .A2(_04299_),
    .B(_04307_),
    .ZN(_01076_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08901_ (.A1(_02612_),
    .A2(_04197_),
    .ZN(_04308_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08902_ (.I(_04308_),
    .Z(_04309_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08903_ (.A1(\u_cpu.rf_ram.memory[96][0] ),
    .A2(_04309_),
    .ZN(_04310_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08904_ (.A1(_04280_),
    .A2(_04309_),
    .B(_04310_),
    .ZN(_01077_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08905_ (.A1(\u_cpu.rf_ram.memory[96][1] ),
    .A2(_04309_),
    .ZN(_04311_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08906_ (.A1(_04284_),
    .A2(_04309_),
    .B(_04311_),
    .ZN(_01078_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08907_ (.A1(\u_cpu.rf_ram.memory[96][2] ),
    .A2(_04309_),
    .ZN(_04312_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08908_ (.A1(_04286_),
    .A2(_04309_),
    .B(_04312_),
    .ZN(_01079_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08909_ (.A1(\u_cpu.rf_ram.memory[96][3] ),
    .A2(_04309_),
    .ZN(_04313_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08910_ (.A1(_04288_),
    .A2(_04309_),
    .B(_04313_),
    .ZN(_01080_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08911_ (.A1(\u_cpu.rf_ram.memory[96][4] ),
    .A2(_04309_),
    .ZN(_04314_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08912_ (.A1(_04290_),
    .A2(_04309_),
    .B(_04314_),
    .ZN(_01081_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08913_ (.A1(\u_cpu.rf_ram.memory[96][5] ),
    .A2(_04309_),
    .ZN(_04315_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08914_ (.A1(_04292_),
    .A2(_04309_),
    .B(_04315_),
    .ZN(_01082_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08915_ (.A1(\u_cpu.rf_ram.memory[96][6] ),
    .A2(_04309_),
    .ZN(_04316_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08916_ (.A1(_04294_),
    .A2(_04309_),
    .B(_04316_),
    .ZN(_01083_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08917_ (.A1(\u_cpu.rf_ram.memory[96][7] ),
    .A2(_04309_),
    .ZN(_04317_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08918_ (.A1(_04296_),
    .A2(_04309_),
    .B(_04317_),
    .ZN(_01084_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08919_ (.A1(\u_cpu.cpu.bufreg.i_sh_signed ),
    .A2(_03798_),
    .ZN(_04318_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08920_ (.A1(_03991_),
    .A2(_04318_),
    .ZN(_01085_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08921_ (.A1(\u_arbiter.i_wb_cpu_ack ),
    .A2(\u_arbiter.o_wb_cpu_adr[1] ),
    .ZN(_04319_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08922_ (.A1(_01437_),
    .A2(_04319_),
    .Z(_04320_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08923_ (.A1(_01428_),
    .A2(_04320_),
    .ZN(_01086_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08924_ (.A1(_02528_),
    .A2(_02671_),
    .ZN(_04321_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08925_ (.I(_04321_),
    .Z(_04322_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08926_ (.A1(\u_cpu.rf_ram.memory[28][0] ),
    .A2(_04322_),
    .ZN(_04323_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08927_ (.A1(_04280_),
    .A2(_04322_),
    .B(_04323_),
    .ZN(_01087_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08928_ (.A1(\u_cpu.rf_ram.memory[28][1] ),
    .A2(_04322_),
    .ZN(_04324_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08929_ (.A1(_04284_),
    .A2(_04322_),
    .B(_04324_),
    .ZN(_01088_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08930_ (.A1(\u_cpu.rf_ram.memory[28][2] ),
    .A2(_04322_),
    .ZN(_04325_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08931_ (.A1(_04286_),
    .A2(_04322_),
    .B(_04325_),
    .ZN(_01089_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08932_ (.A1(\u_cpu.rf_ram.memory[28][3] ),
    .A2(_04322_),
    .ZN(_04326_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08933_ (.A1(_04288_),
    .A2(_04322_),
    .B(_04326_),
    .ZN(_01090_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08934_ (.A1(\u_cpu.rf_ram.memory[28][4] ),
    .A2(_04322_),
    .ZN(_04327_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08935_ (.A1(_04290_),
    .A2(_04322_),
    .B(_04327_),
    .ZN(_01091_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08936_ (.A1(\u_cpu.rf_ram.memory[28][5] ),
    .A2(_04322_),
    .ZN(_04328_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08937_ (.A1(_04292_),
    .A2(_04322_),
    .B(_04328_),
    .ZN(_01092_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08938_ (.A1(\u_cpu.rf_ram.memory[28][6] ),
    .A2(_04322_),
    .ZN(_04329_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08939_ (.A1(_04294_),
    .A2(_04322_),
    .B(_04329_),
    .ZN(_01093_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08940_ (.A1(\u_cpu.rf_ram.memory[28][7] ),
    .A2(_04322_),
    .ZN(_04330_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08941_ (.A1(_04296_),
    .A2(_04322_),
    .B(_04330_),
    .ZN(_01094_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08942_ (.I(_02766_),
    .Z(_04331_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08943_ (.I0(\u_arbiter.i_wb_cpu_rdt[16] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[0] ),
    .S(_04331_),
    .Z(_04332_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08944_ (.I(_04332_),
    .Z(_01095_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08945_ (.I0(\u_arbiter.i_wb_cpu_rdt[17] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[1] ),
    .S(_04331_),
    .Z(_04333_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08946_ (.I(_04333_),
    .Z(_01096_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08947_ (.I0(\u_arbiter.i_wb_cpu_rdt[18] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[2] ),
    .S(_04331_),
    .Z(_04334_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08948_ (.I(_04334_),
    .Z(_01097_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08949_ (.I0(\u_arbiter.i_wb_cpu_rdt[19] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[3] ),
    .S(_04331_),
    .Z(_04335_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08950_ (.I(_04335_),
    .Z(_01098_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08951_ (.I0(\u_arbiter.i_wb_cpu_rdt[20] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[4] ),
    .S(_04331_),
    .Z(_04336_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08952_ (.I(_04336_),
    .Z(_01099_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08953_ (.I0(\u_arbiter.i_wb_cpu_rdt[21] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[5] ),
    .S(_04331_),
    .Z(_04337_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08954_ (.I(_04337_),
    .Z(_01100_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08955_ (.I0(\u_arbiter.i_wb_cpu_rdt[22] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[6] ),
    .S(_04331_),
    .Z(_04338_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08956_ (.I(_04338_),
    .Z(_01101_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08957_ (.I0(\u_arbiter.i_wb_cpu_rdt[23] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[7] ),
    .S(_04331_),
    .Z(_04339_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08958_ (.I(_04339_),
    .Z(_01102_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08959_ (.I0(\u_arbiter.i_wb_cpu_rdt[24] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[8] ),
    .S(_04331_),
    .Z(_04340_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08960_ (.I(_04340_),
    .Z(_01103_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08961_ (.I0(\u_arbiter.i_wb_cpu_rdt[25] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[9] ),
    .S(_04331_),
    .Z(_04341_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08962_ (.I(_04341_),
    .Z(_01104_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08963_ (.I0(\u_arbiter.i_wb_cpu_rdt[26] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[10] ),
    .S(_04331_),
    .Z(_04342_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08964_ (.I(_04342_),
    .Z(_01105_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08965_ (.I0(\u_arbiter.i_wb_cpu_rdt[27] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[11] ),
    .S(_04331_),
    .Z(_04343_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08966_ (.I(_04343_),
    .Z(_01106_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08967_ (.I0(\u_arbiter.i_wb_cpu_rdt[28] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[12] ),
    .S(_04331_),
    .Z(_04344_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08968_ (.I(_04344_),
    .Z(_01107_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08969_ (.I0(\u_arbiter.i_wb_cpu_rdt[29] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[13] ),
    .S(_04331_),
    .Z(_04345_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08970_ (.I(_04345_),
    .Z(_01108_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08971_ (.I0(\u_arbiter.i_wb_cpu_rdt[30] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[14] ),
    .S(_04331_),
    .Z(_04346_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08972_ (.I(_04346_),
    .Z(_01109_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08973_ (.I0(\u_arbiter.i_wb_cpu_rdt[31] ),
    .I1(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[15] ),
    .S(_04331_),
    .Z(_04347_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08974_ (.I(_04347_),
    .Z(_01110_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08975_ (.A1(_02524_),
    .A2(_04197_),
    .ZN(_04348_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08976_ (.I(_04348_),
    .Z(_04349_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08977_ (.A1(\u_cpu.rf_ram.memory[101][0] ),
    .A2(_04349_),
    .ZN(_04350_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08978_ (.A1(_04280_),
    .A2(_04349_),
    .B(_04350_),
    .ZN(_01111_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08979_ (.A1(\u_cpu.rf_ram.memory[101][1] ),
    .A2(_04349_),
    .ZN(_04351_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08980_ (.A1(_04284_),
    .A2(_04349_),
    .B(_04351_),
    .ZN(_01112_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08981_ (.A1(\u_cpu.rf_ram.memory[101][2] ),
    .A2(_04349_),
    .ZN(_04352_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08982_ (.A1(_04286_),
    .A2(_04349_),
    .B(_04352_),
    .ZN(_01113_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08983_ (.A1(\u_cpu.rf_ram.memory[101][3] ),
    .A2(_04349_),
    .ZN(_04353_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08984_ (.A1(_04288_),
    .A2(_04349_),
    .B(_04353_),
    .ZN(_01114_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08985_ (.A1(\u_cpu.rf_ram.memory[101][4] ),
    .A2(_04349_),
    .ZN(_04354_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08986_ (.A1(_04290_),
    .A2(_04349_),
    .B(_04354_),
    .ZN(_01115_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08987_ (.A1(\u_cpu.rf_ram.memory[101][5] ),
    .A2(_04349_),
    .ZN(_04355_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08988_ (.A1(_04292_),
    .A2(_04349_),
    .B(_04355_),
    .ZN(_01116_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08989_ (.A1(\u_cpu.rf_ram.memory[101][6] ),
    .A2(_04349_),
    .ZN(_04356_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08990_ (.A1(_04294_),
    .A2(_04349_),
    .B(_04356_),
    .ZN(_01117_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08991_ (.A1(\u_cpu.rf_ram.memory[101][7] ),
    .A2(_04349_),
    .ZN(_04357_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08992_ (.A1(_04296_),
    .A2(_04349_),
    .B(_04357_),
    .ZN(_01118_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08993_ (.A1(_02893_),
    .A2(_04197_),
    .ZN(_04358_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08994_ (.I(_04358_),
    .Z(_04359_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08995_ (.A1(\u_cpu.rf_ram.memory[102][0] ),
    .A2(_04359_),
    .ZN(_04360_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08996_ (.A1(_04280_),
    .A2(_04359_),
    .B(_04360_),
    .ZN(_01119_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08997_ (.A1(\u_cpu.rf_ram.memory[102][1] ),
    .A2(_04359_),
    .ZN(_04361_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08998_ (.A1(_04284_),
    .A2(_04359_),
    .B(_04361_),
    .ZN(_01120_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08999_ (.A1(\u_cpu.rf_ram.memory[102][2] ),
    .A2(_04359_),
    .ZN(_04362_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09000_ (.A1(_04286_),
    .A2(_04359_),
    .B(_04362_),
    .ZN(_01121_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09001_ (.A1(\u_cpu.rf_ram.memory[102][3] ),
    .A2(_04359_),
    .ZN(_04363_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09002_ (.A1(_04288_),
    .A2(_04359_),
    .B(_04363_),
    .ZN(_01122_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09003_ (.A1(\u_cpu.rf_ram.memory[102][4] ),
    .A2(_04359_),
    .ZN(_04364_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09004_ (.A1(_04290_),
    .A2(_04359_),
    .B(_04364_),
    .ZN(_01123_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09005_ (.A1(\u_cpu.rf_ram.memory[102][5] ),
    .A2(_04359_),
    .ZN(_04365_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09006_ (.A1(_04292_),
    .A2(_04359_),
    .B(_04365_),
    .ZN(_01124_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09007_ (.A1(\u_cpu.rf_ram.memory[102][6] ),
    .A2(_04359_),
    .ZN(_04366_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09008_ (.A1(_04294_),
    .A2(_04359_),
    .B(_04366_),
    .ZN(_01125_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09009_ (.A1(\u_cpu.rf_ram.memory[102][7] ),
    .A2(_04359_),
    .ZN(_04367_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09010_ (.A1(_04296_),
    .A2(_04359_),
    .B(_04367_),
    .ZN(_01126_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09011_ (.A1(_02602_),
    .A2(_04197_),
    .ZN(_04368_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09012_ (.I(_04368_),
    .Z(_04369_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09013_ (.A1(\u_cpu.rf_ram.memory[103][0] ),
    .A2(_04369_),
    .ZN(_04370_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09014_ (.A1(_04280_),
    .A2(_04369_),
    .B(_04370_),
    .ZN(_01127_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09015_ (.A1(\u_cpu.rf_ram.memory[103][1] ),
    .A2(_04369_),
    .ZN(_04371_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09016_ (.A1(_04284_),
    .A2(_04369_),
    .B(_04371_),
    .ZN(_01128_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09017_ (.A1(\u_cpu.rf_ram.memory[103][2] ),
    .A2(_04369_),
    .ZN(_04372_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09018_ (.A1(_04286_),
    .A2(_04369_),
    .B(_04372_),
    .ZN(_01129_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09019_ (.A1(\u_cpu.rf_ram.memory[103][3] ),
    .A2(_04369_),
    .ZN(_04373_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09020_ (.A1(_04288_),
    .A2(_04369_),
    .B(_04373_),
    .ZN(_01130_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09021_ (.A1(\u_cpu.rf_ram.memory[103][4] ),
    .A2(_04369_),
    .ZN(_04374_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09022_ (.A1(_04290_),
    .A2(_04369_),
    .B(_04374_),
    .ZN(_01131_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09023_ (.A1(\u_cpu.rf_ram.memory[103][5] ),
    .A2(_04369_),
    .ZN(_04375_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09024_ (.A1(_04292_),
    .A2(_04369_),
    .B(_04375_),
    .ZN(_01132_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09025_ (.A1(\u_cpu.rf_ram.memory[103][6] ),
    .A2(_04369_),
    .ZN(_04376_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09026_ (.A1(_04294_),
    .A2(_04369_),
    .B(_04376_),
    .ZN(_01133_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09027_ (.A1(\u_cpu.rf_ram.memory[103][7] ),
    .A2(_04369_),
    .ZN(_04377_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09028_ (.A1(_04296_),
    .A2(_04369_),
    .B(_04377_),
    .ZN(_01134_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09029_ (.A1(_02810_),
    .A2(_04197_),
    .ZN(_04378_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09030_ (.I(_04378_),
    .Z(_04379_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09031_ (.A1(\u_cpu.rf_ram.memory[104][0] ),
    .A2(_04379_),
    .ZN(_04380_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09032_ (.A1(_04280_),
    .A2(_04379_),
    .B(_04380_),
    .ZN(_01135_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09033_ (.A1(\u_cpu.rf_ram.memory[104][1] ),
    .A2(_04379_),
    .ZN(_04381_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09034_ (.A1(_04284_),
    .A2(_04379_),
    .B(_04381_),
    .ZN(_01136_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09035_ (.A1(\u_cpu.rf_ram.memory[104][2] ),
    .A2(_04379_),
    .ZN(_04382_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09036_ (.A1(_04286_),
    .A2(_04379_),
    .B(_04382_),
    .ZN(_01137_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09037_ (.A1(\u_cpu.rf_ram.memory[104][3] ),
    .A2(_04379_),
    .ZN(_04383_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09038_ (.A1(_04288_),
    .A2(_04379_),
    .B(_04383_),
    .ZN(_01138_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09039_ (.A1(\u_cpu.rf_ram.memory[104][4] ),
    .A2(_04379_),
    .ZN(_04384_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09040_ (.A1(_04290_),
    .A2(_04379_),
    .B(_04384_),
    .ZN(_01139_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09041_ (.A1(\u_cpu.rf_ram.memory[104][5] ),
    .A2(_04379_),
    .ZN(_04385_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09042_ (.A1(_04292_),
    .A2(_04379_),
    .B(_04385_),
    .ZN(_01140_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09043_ (.A1(\u_cpu.rf_ram.memory[104][6] ),
    .A2(_04379_),
    .ZN(_04386_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09044_ (.A1(_04294_),
    .A2(_04379_),
    .B(_04386_),
    .ZN(_01141_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09045_ (.A1(\u_cpu.rf_ram.memory[104][7] ),
    .A2(_04379_),
    .ZN(_04387_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09046_ (.A1(_04296_),
    .A2(_04379_),
    .B(_04387_),
    .ZN(_01142_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09047_ (.A1(_02682_),
    .A2(_04197_),
    .ZN(_04388_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09048_ (.I(_04388_),
    .Z(_04389_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09049_ (.A1(\u_cpu.rf_ram.memory[99][0] ),
    .A2(_04389_),
    .ZN(_04390_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09050_ (.A1(_04280_),
    .A2(_04389_),
    .B(_04390_),
    .ZN(_01143_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09051_ (.A1(\u_cpu.rf_ram.memory[99][1] ),
    .A2(_04389_),
    .ZN(_04391_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09052_ (.A1(_04284_),
    .A2(_04389_),
    .B(_04391_),
    .ZN(_01144_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09053_ (.A1(\u_cpu.rf_ram.memory[99][2] ),
    .A2(_04389_),
    .ZN(_04392_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09054_ (.A1(_04286_),
    .A2(_04389_),
    .B(_04392_),
    .ZN(_01145_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09055_ (.A1(\u_cpu.rf_ram.memory[99][3] ),
    .A2(_04389_),
    .ZN(_04393_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09056_ (.A1(_04288_),
    .A2(_04389_),
    .B(_04393_),
    .ZN(_01146_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09057_ (.A1(\u_cpu.rf_ram.memory[99][4] ),
    .A2(_04389_),
    .ZN(_04394_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09058_ (.A1(_04290_),
    .A2(_04389_),
    .B(_04394_),
    .ZN(_01147_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09059_ (.A1(\u_cpu.rf_ram.memory[99][5] ),
    .A2(_04389_),
    .ZN(_04395_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09060_ (.A1(_04292_),
    .A2(_04389_),
    .B(_04395_),
    .ZN(_01148_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09061_ (.A1(\u_cpu.rf_ram.memory[99][6] ),
    .A2(_04389_),
    .ZN(_04396_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09062_ (.A1(_04294_),
    .A2(_04389_),
    .B(_04396_),
    .ZN(_01149_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09063_ (.A1(\u_cpu.rf_ram.memory[99][7] ),
    .A2(_04389_),
    .ZN(_04397_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09064_ (.A1(_04296_),
    .A2(_04389_),
    .B(_04397_),
    .ZN(_01150_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09065_ (.A1(_02626_),
    .A2(_02727_),
    .ZN(_04398_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09066_ (.I(_04398_),
    .Z(_04399_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09067_ (.A1(\u_cpu.rf_ram.memory[79][0] ),
    .A2(_04399_),
    .ZN(_04400_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09068_ (.A1(_04280_),
    .A2(_04399_),
    .B(_04400_),
    .ZN(_01151_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09069_ (.A1(\u_cpu.rf_ram.memory[79][1] ),
    .A2(_04399_),
    .ZN(_04401_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09070_ (.A1(_04284_),
    .A2(_04399_),
    .B(_04401_),
    .ZN(_01152_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09071_ (.A1(\u_cpu.rf_ram.memory[79][2] ),
    .A2(_04399_),
    .ZN(_04402_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09072_ (.A1(_04286_),
    .A2(_04399_),
    .B(_04402_),
    .ZN(_01153_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09073_ (.A1(\u_cpu.rf_ram.memory[79][3] ),
    .A2(_04399_),
    .ZN(_04403_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09074_ (.A1(_04288_),
    .A2(_04399_),
    .B(_04403_),
    .ZN(_01154_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09075_ (.A1(\u_cpu.rf_ram.memory[79][4] ),
    .A2(_04399_),
    .ZN(_04404_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09076_ (.A1(_04290_),
    .A2(_04399_),
    .B(_04404_),
    .ZN(_01155_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09077_ (.A1(\u_cpu.rf_ram.memory[79][5] ),
    .A2(_04399_),
    .ZN(_04405_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09078_ (.A1(_04292_),
    .A2(_04399_),
    .B(_04405_),
    .ZN(_01156_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09079_ (.A1(\u_cpu.rf_ram.memory[79][6] ),
    .A2(_04399_),
    .ZN(_04406_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09080_ (.A1(_04294_),
    .A2(_04399_),
    .B(_04406_),
    .ZN(_01157_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09081_ (.A1(\u_cpu.rf_ram.memory[79][7] ),
    .A2(_04399_),
    .ZN(_04407_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09082_ (.A1(_04296_),
    .A2(_04399_),
    .B(_04407_),
    .ZN(_01158_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09083_ (.A1(_02695_),
    .A2(_04197_),
    .ZN(_04408_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09084_ (.I(_04408_),
    .Z(_04409_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09085_ (.A1(\u_cpu.rf_ram.memory[105][0] ),
    .A2(_04409_),
    .ZN(_04410_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09086_ (.A1(_04280_),
    .A2(_04409_),
    .B(_04410_),
    .ZN(_01159_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09087_ (.A1(\u_cpu.rf_ram.memory[105][1] ),
    .A2(_04409_),
    .ZN(_04411_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09088_ (.A1(_04284_),
    .A2(_04409_),
    .B(_04411_),
    .ZN(_01160_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09089_ (.A1(\u_cpu.rf_ram.memory[105][2] ),
    .A2(_04409_),
    .ZN(_04412_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09090_ (.A1(_04286_),
    .A2(_04409_),
    .B(_04412_),
    .ZN(_01161_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09091_ (.A1(\u_cpu.rf_ram.memory[105][3] ),
    .A2(_04409_),
    .ZN(_04413_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09092_ (.A1(_04288_),
    .A2(_04409_),
    .B(_04413_),
    .ZN(_01162_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09093_ (.A1(\u_cpu.rf_ram.memory[105][4] ),
    .A2(_04409_),
    .ZN(_04414_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09094_ (.A1(_04290_),
    .A2(_04409_),
    .B(_04414_),
    .ZN(_01163_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09095_ (.A1(\u_cpu.rf_ram.memory[105][5] ),
    .A2(_04409_),
    .ZN(_04415_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09096_ (.A1(_04292_),
    .A2(_04409_),
    .B(_04415_),
    .ZN(_01164_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09097_ (.A1(\u_cpu.rf_ram.memory[105][6] ),
    .A2(_04409_),
    .ZN(_04416_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09098_ (.A1(_04294_),
    .A2(_04409_),
    .B(_04416_),
    .ZN(_01165_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09099_ (.A1(\u_cpu.rf_ram.memory[105][7] ),
    .A2(_04409_),
    .ZN(_04417_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09100_ (.A1(_04296_),
    .A2(_04409_),
    .B(_04417_),
    .ZN(_01166_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09101_ (.A1(_02638_),
    .A2(_04197_),
    .ZN(_04418_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09102_ (.I(_04418_),
    .Z(_04419_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09103_ (.A1(\u_cpu.rf_ram.memory[106][0] ),
    .A2(_04419_),
    .ZN(_04420_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09104_ (.A1(_04280_),
    .A2(_04419_),
    .B(_04420_),
    .ZN(_01167_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09105_ (.A1(\u_cpu.rf_ram.memory[106][1] ),
    .A2(_04419_),
    .ZN(_04421_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09106_ (.A1(_04284_),
    .A2(_04419_),
    .B(_04421_),
    .ZN(_01168_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09107_ (.A1(\u_cpu.rf_ram.memory[106][2] ),
    .A2(_04419_),
    .ZN(_04422_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09108_ (.A1(_04286_),
    .A2(_04419_),
    .B(_04422_),
    .ZN(_01169_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09109_ (.A1(\u_cpu.rf_ram.memory[106][3] ),
    .A2(_04419_),
    .ZN(_04423_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09110_ (.A1(_04288_),
    .A2(_04419_),
    .B(_04423_),
    .ZN(_01170_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09111_ (.A1(\u_cpu.rf_ram.memory[106][4] ),
    .A2(_04419_),
    .ZN(_04424_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09112_ (.A1(_04290_),
    .A2(_04419_),
    .B(_04424_),
    .ZN(_01171_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09113_ (.A1(\u_cpu.rf_ram.memory[106][5] ),
    .A2(_04419_),
    .ZN(_04425_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09114_ (.A1(_04292_),
    .A2(_04419_),
    .B(_04425_),
    .ZN(_01172_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09115_ (.A1(\u_cpu.rf_ram.memory[106][6] ),
    .A2(_04419_),
    .ZN(_04426_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09116_ (.A1(_04294_),
    .A2(_04419_),
    .B(_04426_),
    .ZN(_01173_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09117_ (.A1(\u_cpu.rf_ram.memory[106][7] ),
    .A2(_04419_),
    .ZN(_04427_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09118_ (.A1(_04296_),
    .A2(_04419_),
    .B(_04427_),
    .ZN(_01174_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09119_ (.A1(_02706_),
    .A2(_04197_),
    .ZN(_04428_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09120_ (.I(_04428_),
    .Z(_04429_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09121_ (.A1(\u_cpu.rf_ram.memory[107][0] ),
    .A2(_04429_),
    .ZN(_04430_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09122_ (.A1(_04280_),
    .A2(_04429_),
    .B(_04430_),
    .ZN(_01175_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09123_ (.A1(\u_cpu.rf_ram.memory[107][1] ),
    .A2(_04429_),
    .ZN(_04431_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09124_ (.A1(_04284_),
    .A2(_04429_),
    .B(_04431_),
    .ZN(_01176_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09125_ (.A1(\u_cpu.rf_ram.memory[107][2] ),
    .A2(_04429_),
    .ZN(_04432_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09126_ (.A1(_04286_),
    .A2(_04429_),
    .B(_04432_),
    .ZN(_01177_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09127_ (.A1(\u_cpu.rf_ram.memory[107][3] ),
    .A2(_04429_),
    .ZN(_04433_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09128_ (.A1(_04288_),
    .A2(_04429_),
    .B(_04433_),
    .ZN(_01178_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09129_ (.A1(\u_cpu.rf_ram.memory[107][4] ),
    .A2(_04429_),
    .ZN(_04434_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09130_ (.A1(_04290_),
    .A2(_04429_),
    .B(_04434_),
    .ZN(_01179_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09131_ (.A1(\u_cpu.rf_ram.memory[107][5] ),
    .A2(_04429_),
    .ZN(_04435_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09132_ (.A1(_04292_),
    .A2(_04429_),
    .B(_04435_),
    .ZN(_01180_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09133_ (.A1(\u_cpu.rf_ram.memory[107][6] ),
    .A2(_04429_),
    .ZN(_04436_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09134_ (.A1(_04294_),
    .A2(_04429_),
    .B(_04436_),
    .ZN(_01181_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09135_ (.A1(\u_cpu.rf_ram.memory[107][7] ),
    .A2(_04429_),
    .ZN(_04437_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09136_ (.A1(_04296_),
    .A2(_04429_),
    .B(_04437_),
    .ZN(_01182_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09137_ (.A1(_02475_),
    .A2(_02682_),
    .ZN(_04438_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09138_ (.I(_04438_),
    .Z(_04439_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09139_ (.A1(\u_cpu.rf_ram.memory[83][0] ),
    .A2(_04439_),
    .ZN(_04440_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09140_ (.A1(_04280_),
    .A2(_04439_),
    .B(_04440_),
    .ZN(_01183_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09141_ (.A1(\u_cpu.rf_ram.memory[83][1] ),
    .A2(_04439_),
    .ZN(_04441_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09142_ (.A1(_04284_),
    .A2(_04439_),
    .B(_04441_),
    .ZN(_01184_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09143_ (.A1(\u_cpu.rf_ram.memory[83][2] ),
    .A2(_04439_),
    .ZN(_04442_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09144_ (.A1(_04286_),
    .A2(_04439_),
    .B(_04442_),
    .ZN(_01185_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09145_ (.A1(\u_cpu.rf_ram.memory[83][3] ),
    .A2(_04439_),
    .ZN(_04443_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09146_ (.A1(_04288_),
    .A2(_04439_),
    .B(_04443_),
    .ZN(_01186_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09147_ (.A1(\u_cpu.rf_ram.memory[83][4] ),
    .A2(_04439_),
    .ZN(_04444_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09148_ (.A1(_04290_),
    .A2(_04439_),
    .B(_04444_),
    .ZN(_01187_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09149_ (.A1(\u_cpu.rf_ram.memory[83][5] ),
    .A2(_04439_),
    .ZN(_04445_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09150_ (.A1(_04292_),
    .A2(_04439_),
    .B(_04445_),
    .ZN(_01188_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09151_ (.A1(\u_cpu.rf_ram.memory[83][6] ),
    .A2(_04439_),
    .ZN(_04446_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09152_ (.A1(_04294_),
    .A2(_04439_),
    .B(_04446_),
    .ZN(_01189_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09153_ (.A1(\u_cpu.rf_ram.memory[83][7] ),
    .A2(_04439_),
    .ZN(_04447_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09154_ (.A1(_04296_),
    .A2(_04439_),
    .B(_04447_),
    .ZN(_01190_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09155_ (.A1(_02671_),
    .A2(_04197_),
    .ZN(_04448_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09156_ (.I(_04448_),
    .Z(_04449_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09157_ (.A1(\u_cpu.rf_ram.memory[108][0] ),
    .A2(_04449_),
    .ZN(_04450_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09158_ (.A1(_04280_),
    .A2(_04449_),
    .B(_04450_),
    .ZN(_01191_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09159_ (.A1(\u_cpu.rf_ram.memory[108][1] ),
    .A2(_04449_),
    .ZN(_04451_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09160_ (.A1(_04284_),
    .A2(_04449_),
    .B(_04451_),
    .ZN(_01192_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09161_ (.A1(\u_cpu.rf_ram.memory[108][2] ),
    .A2(_04449_),
    .ZN(_04452_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09162_ (.A1(_04286_),
    .A2(_04449_),
    .B(_04452_),
    .ZN(_01193_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09163_ (.A1(\u_cpu.rf_ram.memory[108][3] ),
    .A2(_04449_),
    .ZN(_04453_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09164_ (.A1(_04288_),
    .A2(_04449_),
    .B(_04453_),
    .ZN(_01194_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09165_ (.A1(\u_cpu.rf_ram.memory[108][4] ),
    .A2(_04449_),
    .ZN(_04454_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09166_ (.A1(_04290_),
    .A2(_04449_),
    .B(_04454_),
    .ZN(_01195_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09167_ (.A1(\u_cpu.rf_ram.memory[108][5] ),
    .A2(_04449_),
    .ZN(_04455_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09168_ (.A1(_04292_),
    .A2(_04449_),
    .B(_04455_),
    .ZN(_01196_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09169_ (.A1(\u_cpu.rf_ram.memory[108][6] ),
    .A2(_04449_),
    .ZN(_04456_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09170_ (.A1(_04294_),
    .A2(_04449_),
    .B(_04456_),
    .ZN(_01197_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09171_ (.A1(\u_cpu.rf_ram.memory[108][7] ),
    .A2(_04449_),
    .ZN(_04457_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09172_ (.A1(_04296_),
    .A2(_04449_),
    .B(_04457_),
    .ZN(_01198_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09173_ (.A1(_02524_),
    .A2(_02626_),
    .ZN(_04458_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09174_ (.I(_04458_),
    .Z(_04459_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09175_ (.A1(\u_cpu.rf_ram.memory[69][0] ),
    .A2(_04459_),
    .ZN(_04460_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09176_ (.A1(_04280_),
    .A2(_04459_),
    .B(_04460_),
    .ZN(_01199_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09177_ (.A1(\u_cpu.rf_ram.memory[69][1] ),
    .A2(_04459_),
    .ZN(_04461_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09178_ (.A1(_04284_),
    .A2(_04459_),
    .B(_04461_),
    .ZN(_01200_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09179_ (.A1(\u_cpu.rf_ram.memory[69][2] ),
    .A2(_04459_),
    .ZN(_04462_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09180_ (.A1(_04286_),
    .A2(_04459_),
    .B(_04462_),
    .ZN(_01201_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09181_ (.A1(\u_cpu.rf_ram.memory[69][3] ),
    .A2(_04459_),
    .ZN(_04463_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09182_ (.A1(_04288_),
    .A2(_04459_),
    .B(_04463_),
    .ZN(_01202_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09183_ (.A1(\u_cpu.rf_ram.memory[69][4] ),
    .A2(_04459_),
    .ZN(_04464_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09184_ (.A1(_04290_),
    .A2(_04459_),
    .B(_04464_),
    .ZN(_01203_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09185_ (.A1(\u_cpu.rf_ram.memory[69][5] ),
    .A2(_04459_),
    .ZN(_04465_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09186_ (.A1(_04292_),
    .A2(_04459_),
    .B(_04465_),
    .ZN(_01204_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09187_ (.A1(\u_cpu.rf_ram.memory[69][6] ),
    .A2(_04459_),
    .ZN(_04466_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09188_ (.A1(_04294_),
    .A2(_04459_),
    .B(_04466_),
    .ZN(_01205_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09189_ (.A1(\u_cpu.rf_ram.memory[69][7] ),
    .A2(_04459_),
    .ZN(_04467_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09190_ (.A1(_04296_),
    .A2(_04459_),
    .B(_04467_),
    .ZN(_01206_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09191_ (.I(_02481_),
    .Z(_04468_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09192_ (.A1(_02475_),
    .A2(_02561_),
    .ZN(_04469_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09193_ (.I(_04469_),
    .Z(_04470_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09194_ (.A1(\u_cpu.rf_ram.memory[84][0] ),
    .A2(_04470_),
    .ZN(_04471_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09195_ (.A1(_04468_),
    .A2(_04470_),
    .B(_04471_),
    .ZN(_01207_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09196_ (.I(_02486_),
    .Z(_04472_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09197_ (.A1(\u_cpu.rf_ram.memory[84][1] ),
    .A2(_04470_),
    .ZN(_04473_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09198_ (.A1(_04472_),
    .A2(_04470_),
    .B(_04473_),
    .ZN(_01208_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09199_ (.I(_02491_),
    .Z(_04474_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09200_ (.A1(\u_cpu.rf_ram.memory[84][2] ),
    .A2(_04470_),
    .ZN(_04475_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09201_ (.A1(_04474_),
    .A2(_04470_),
    .B(_04475_),
    .ZN(_01209_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09202_ (.I(_02496_),
    .Z(_04476_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09203_ (.A1(\u_cpu.rf_ram.memory[84][3] ),
    .A2(_04470_),
    .ZN(_04477_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09204_ (.A1(_04476_),
    .A2(_04470_),
    .B(_04477_),
    .ZN(_01210_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09205_ (.I(_02501_),
    .Z(_04478_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09206_ (.A1(\u_cpu.rf_ram.memory[84][4] ),
    .A2(_04470_),
    .ZN(_04479_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09207_ (.A1(_04478_),
    .A2(_04470_),
    .B(_04479_),
    .ZN(_01211_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09208_ (.I(_02506_),
    .Z(_04480_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09209_ (.A1(\u_cpu.rf_ram.memory[84][5] ),
    .A2(_04470_),
    .ZN(_04481_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09210_ (.A1(_04480_),
    .A2(_04470_),
    .B(_04481_),
    .ZN(_01212_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09211_ (.I(_02511_),
    .Z(_04482_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09212_ (.A1(\u_cpu.rf_ram.memory[84][6] ),
    .A2(_04470_),
    .ZN(_04483_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09213_ (.A1(_04482_),
    .A2(_04470_),
    .B(_04483_),
    .ZN(_01213_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09214_ (.I(_02516_),
    .Z(_04484_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09215_ (.A1(\u_cpu.rf_ram.memory[84][7] ),
    .A2(_04470_),
    .ZN(_04485_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09216_ (.A1(_04484_),
    .A2(_04470_),
    .B(_04485_),
    .ZN(_01214_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09217_ (.A1(_02684_),
    .A2(_02706_),
    .ZN(_04486_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09218_ (.I(_04486_),
    .Z(_04487_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09219_ (.A1(\u_cpu.rf_ram.memory[59][0] ),
    .A2(_04487_),
    .ZN(_04488_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09220_ (.A1(_04468_),
    .A2(_04487_),
    .B(_04488_),
    .ZN(_01215_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09221_ (.A1(\u_cpu.rf_ram.memory[59][1] ),
    .A2(_04487_),
    .ZN(_04489_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09222_ (.A1(_04472_),
    .A2(_04487_),
    .B(_04489_),
    .ZN(_01216_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09223_ (.A1(\u_cpu.rf_ram.memory[59][2] ),
    .A2(_04487_),
    .ZN(_04490_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09224_ (.A1(_04474_),
    .A2(_04487_),
    .B(_04490_),
    .ZN(_01217_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09225_ (.A1(\u_cpu.rf_ram.memory[59][3] ),
    .A2(_04487_),
    .ZN(_04491_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09226_ (.A1(_04476_),
    .A2(_04487_),
    .B(_04491_),
    .ZN(_01218_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09227_ (.A1(\u_cpu.rf_ram.memory[59][4] ),
    .A2(_04487_),
    .ZN(_04492_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09228_ (.A1(_04478_),
    .A2(_04487_),
    .B(_04492_),
    .ZN(_01219_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09229_ (.A1(\u_cpu.rf_ram.memory[59][5] ),
    .A2(_04487_),
    .ZN(_04493_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09230_ (.A1(_04480_),
    .A2(_04487_),
    .B(_04493_),
    .ZN(_01220_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09231_ (.A1(\u_cpu.rf_ram.memory[59][6] ),
    .A2(_04487_),
    .ZN(_04494_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09232_ (.A1(_04482_),
    .A2(_04487_),
    .B(_04494_),
    .ZN(_01221_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09233_ (.A1(\u_cpu.rf_ram.memory[59][7] ),
    .A2(_04487_),
    .ZN(_04495_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09234_ (.A1(_04484_),
    .A2(_04487_),
    .B(_04495_),
    .ZN(_01222_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09235_ (.A1(_02577_),
    .A2(_02638_),
    .ZN(_04496_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09236_ (.I0(_02573_),
    .I1(\u_cpu.rf_ram.memory[10][0] ),
    .S(_04496_),
    .Z(_04497_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09237_ (.I(_04497_),
    .Z(_01223_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09238_ (.I0(_02581_),
    .I1(\u_cpu.rf_ram.memory[10][1] ),
    .S(_04496_),
    .Z(_04498_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09239_ (.I(_04498_),
    .Z(_01224_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09240_ (.I0(_02584_),
    .I1(\u_cpu.rf_ram.memory[10][2] ),
    .S(_04496_),
    .Z(_04499_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09241_ (.I(_04499_),
    .Z(_01225_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09242_ (.I0(_02587_),
    .I1(\u_cpu.rf_ram.memory[10][3] ),
    .S(_04496_),
    .Z(_04500_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09243_ (.I(_04500_),
    .Z(_01226_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09244_ (.I0(_02590_),
    .I1(\u_cpu.rf_ram.memory[10][4] ),
    .S(_04496_),
    .Z(_04501_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09245_ (.I(_04501_),
    .Z(_01227_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09246_ (.I0(_02593_),
    .I1(\u_cpu.rf_ram.memory[10][5] ),
    .S(_04496_),
    .Z(_04502_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09247_ (.I(_04502_),
    .Z(_01228_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09248_ (.I0(_02596_),
    .I1(\u_cpu.rf_ram.memory[10][6] ),
    .S(_04496_),
    .Z(_04503_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09249_ (.I(_04503_),
    .Z(_01229_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09250_ (.I0(_02599_),
    .I1(\u_cpu.rf_ram.memory[10][7] ),
    .S(_04496_),
    .Z(_04504_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09251_ (.I(_04504_),
    .Z(_01230_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09252_ (.A1(_02475_),
    .A2(_02524_),
    .ZN(_04505_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09253_ (.I(_04505_),
    .Z(_04506_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09254_ (.A1(\u_cpu.rf_ram.memory[85][0] ),
    .A2(_04506_),
    .ZN(_04507_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09255_ (.A1(_04468_),
    .A2(_04506_),
    .B(_04507_),
    .ZN(_01231_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09256_ (.A1(\u_cpu.rf_ram.memory[85][1] ),
    .A2(_04506_),
    .ZN(_04508_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09257_ (.A1(_04472_),
    .A2(_04506_),
    .B(_04508_),
    .ZN(_01232_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09258_ (.A1(\u_cpu.rf_ram.memory[85][2] ),
    .A2(_04506_),
    .ZN(_04509_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09259_ (.A1(_04474_),
    .A2(_04506_),
    .B(_04509_),
    .ZN(_01233_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09260_ (.A1(\u_cpu.rf_ram.memory[85][3] ),
    .A2(_04506_),
    .ZN(_04510_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09261_ (.A1(_04476_),
    .A2(_04506_),
    .B(_04510_),
    .ZN(_01234_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09262_ (.A1(\u_cpu.rf_ram.memory[85][4] ),
    .A2(_04506_),
    .ZN(_04511_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09263_ (.A1(_04478_),
    .A2(_04506_),
    .B(_04511_),
    .ZN(_01235_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09264_ (.A1(\u_cpu.rf_ram.memory[85][5] ),
    .A2(_04506_),
    .ZN(_04512_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09265_ (.A1(_04480_),
    .A2(_04506_),
    .B(_04512_),
    .ZN(_01236_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09266_ (.A1(\u_cpu.rf_ram.memory[85][6] ),
    .A2(_04506_),
    .ZN(_04513_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09267_ (.A1(_04482_),
    .A2(_04506_),
    .B(_04513_),
    .ZN(_01237_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09268_ (.A1(\u_cpu.rf_ram.memory[85][7] ),
    .A2(_04506_),
    .ZN(_04514_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09269_ (.A1(_04484_),
    .A2(_04506_),
    .B(_04514_),
    .ZN(_01238_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09270_ (.A1(_02625_),
    .A2(_04197_),
    .ZN(_04515_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09271_ (.I(_04515_),
    .Z(_04516_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09272_ (.A1(\u_cpu.rf_ram.memory[110][0] ),
    .A2(_04516_),
    .ZN(_04517_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09273_ (.A1(_04468_),
    .A2(_04516_),
    .B(_04517_),
    .ZN(_01239_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09274_ (.A1(\u_cpu.rf_ram.memory[110][1] ),
    .A2(_04516_),
    .ZN(_04518_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09275_ (.A1(_04472_),
    .A2(_04516_),
    .B(_04518_),
    .ZN(_01240_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09276_ (.A1(\u_cpu.rf_ram.memory[110][2] ),
    .A2(_04516_),
    .ZN(_04519_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09277_ (.A1(_04474_),
    .A2(_04516_),
    .B(_04519_),
    .ZN(_01241_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09278_ (.A1(\u_cpu.rf_ram.memory[110][3] ),
    .A2(_04516_),
    .ZN(_04520_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09279_ (.A1(_04476_),
    .A2(_04516_),
    .B(_04520_),
    .ZN(_01242_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09280_ (.A1(\u_cpu.rf_ram.memory[110][4] ),
    .A2(_04516_),
    .ZN(_04521_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09281_ (.A1(_04478_),
    .A2(_04516_),
    .B(_04521_),
    .ZN(_01243_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09282_ (.A1(\u_cpu.rf_ram.memory[110][5] ),
    .A2(_04516_),
    .ZN(_04522_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09283_ (.A1(_04480_),
    .A2(_04516_),
    .B(_04522_),
    .ZN(_01244_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09284_ (.A1(\u_cpu.rf_ram.memory[110][6] ),
    .A2(_04516_),
    .ZN(_04523_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09285_ (.A1(_04482_),
    .A2(_04516_),
    .B(_04523_),
    .ZN(_01245_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09286_ (.A1(\u_cpu.rf_ram.memory[110][7] ),
    .A2(_04516_),
    .ZN(_04524_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09287_ (.A1(_04484_),
    .A2(_04516_),
    .B(_04524_),
    .ZN(_01246_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09288_ (.A1(_02475_),
    .A2(_02893_),
    .ZN(_04525_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09289_ (.I(_04525_),
    .Z(_04526_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09290_ (.A1(\u_cpu.rf_ram.memory[86][0] ),
    .A2(_04526_),
    .ZN(_04527_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09291_ (.A1(_04468_),
    .A2(_04526_),
    .B(_04527_),
    .ZN(_01247_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09292_ (.A1(\u_cpu.rf_ram.memory[86][1] ),
    .A2(_04526_),
    .ZN(_04528_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09293_ (.A1(_04472_),
    .A2(_04526_),
    .B(_04528_),
    .ZN(_01248_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09294_ (.A1(\u_cpu.rf_ram.memory[86][2] ),
    .A2(_04526_),
    .ZN(_04529_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09295_ (.A1(_04474_),
    .A2(_04526_),
    .B(_04529_),
    .ZN(_01249_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09296_ (.A1(\u_cpu.rf_ram.memory[86][3] ),
    .A2(_04526_),
    .ZN(_04530_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09297_ (.A1(_04476_),
    .A2(_04526_),
    .B(_04530_),
    .ZN(_01250_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09298_ (.A1(\u_cpu.rf_ram.memory[86][4] ),
    .A2(_04526_),
    .ZN(_04531_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09299_ (.A1(_04478_),
    .A2(_04526_),
    .B(_04531_),
    .ZN(_01251_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09300_ (.A1(\u_cpu.rf_ram.memory[86][5] ),
    .A2(_04526_),
    .ZN(_04532_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09301_ (.A1(_04480_),
    .A2(_04526_),
    .B(_04532_),
    .ZN(_01252_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09302_ (.A1(\u_cpu.rf_ram.memory[86][6] ),
    .A2(_04526_),
    .ZN(_04533_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09303_ (.A1(_04482_),
    .A2(_04526_),
    .B(_04533_),
    .ZN(_01253_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09304_ (.A1(\u_cpu.rf_ram.memory[86][7] ),
    .A2(_04526_),
    .ZN(_04534_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09305_ (.A1(_04484_),
    .A2(_04526_),
    .B(_04534_),
    .ZN(_01254_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09306_ (.A1(_02727_),
    .A2(_04197_),
    .ZN(_04535_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09307_ (.I(_04535_),
    .Z(_04536_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09308_ (.A1(\u_cpu.rf_ram.memory[111][0] ),
    .A2(_04536_),
    .ZN(_04537_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09309_ (.A1(_04468_),
    .A2(_04536_),
    .B(_04537_),
    .ZN(_01255_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09310_ (.A1(\u_cpu.rf_ram.memory[111][1] ),
    .A2(_04536_),
    .ZN(_04538_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09311_ (.A1(_04472_),
    .A2(_04536_),
    .B(_04538_),
    .ZN(_01256_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09312_ (.A1(\u_cpu.rf_ram.memory[111][2] ),
    .A2(_04536_),
    .ZN(_04539_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09313_ (.A1(_04474_),
    .A2(_04536_),
    .B(_04539_),
    .ZN(_01257_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09314_ (.A1(\u_cpu.rf_ram.memory[111][3] ),
    .A2(_04536_),
    .ZN(_04540_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09315_ (.A1(_04476_),
    .A2(_04536_),
    .B(_04540_),
    .ZN(_01258_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09316_ (.A1(\u_cpu.rf_ram.memory[111][4] ),
    .A2(_04536_),
    .ZN(_04541_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09317_ (.A1(_04478_),
    .A2(_04536_),
    .B(_04541_),
    .ZN(_01259_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09318_ (.A1(\u_cpu.rf_ram.memory[111][5] ),
    .A2(_04536_),
    .ZN(_04542_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09319_ (.A1(_04480_),
    .A2(_04536_),
    .B(_04542_),
    .ZN(_01260_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09320_ (.A1(\u_cpu.rf_ram.memory[111][6] ),
    .A2(_04536_),
    .ZN(_04543_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09321_ (.A1(_04482_),
    .A2(_04536_),
    .B(_04543_),
    .ZN(_01261_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09322_ (.A1(\u_cpu.rf_ram.memory[111][7] ),
    .A2(_04536_),
    .ZN(_04544_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09323_ (.A1(_04484_),
    .A2(_04536_),
    .B(_04544_),
    .ZN(_01262_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09324_ (.A1(_02475_),
    .A2(_02602_),
    .ZN(_04545_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09325_ (.I(_04545_),
    .Z(_04546_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09326_ (.A1(\u_cpu.rf_ram.memory[87][0] ),
    .A2(_04546_),
    .ZN(_04547_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09327_ (.A1(_04468_),
    .A2(_04546_),
    .B(_04547_),
    .ZN(_01263_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09328_ (.A1(\u_cpu.rf_ram.memory[87][1] ),
    .A2(_04546_),
    .ZN(_04548_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09329_ (.A1(_04472_),
    .A2(_04546_),
    .B(_04548_),
    .ZN(_01264_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09330_ (.A1(\u_cpu.rf_ram.memory[87][2] ),
    .A2(_04546_),
    .ZN(_04549_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09331_ (.A1(_04474_),
    .A2(_04546_),
    .B(_04549_),
    .ZN(_01265_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09332_ (.A1(\u_cpu.rf_ram.memory[87][3] ),
    .A2(_04546_),
    .ZN(_04550_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09333_ (.A1(_04476_),
    .A2(_04546_),
    .B(_04550_),
    .ZN(_01266_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09334_ (.A1(\u_cpu.rf_ram.memory[87][4] ),
    .A2(_04546_),
    .ZN(_04551_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09335_ (.A1(_04478_),
    .A2(_04546_),
    .B(_04551_),
    .ZN(_01267_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09336_ (.A1(\u_cpu.rf_ram.memory[87][5] ),
    .A2(_04546_),
    .ZN(_04552_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09337_ (.A1(_04480_),
    .A2(_04546_),
    .B(_04552_),
    .ZN(_01268_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09338_ (.A1(\u_cpu.rf_ram.memory[87][6] ),
    .A2(_04546_),
    .ZN(_04553_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09339_ (.A1(_04482_),
    .A2(_04546_),
    .B(_04553_),
    .ZN(_01269_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09340_ (.A1(\u_cpu.rf_ram.memory[87][7] ),
    .A2(_04546_),
    .ZN(_04554_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09341_ (.A1(_04484_),
    .A2(_04546_),
    .B(_04554_),
    .ZN(_01270_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09342_ (.A1(_02475_),
    .A2(_02810_),
    .ZN(_04555_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09343_ (.I(_04555_),
    .Z(_04556_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09344_ (.A1(\u_cpu.rf_ram.memory[88][0] ),
    .A2(_04556_),
    .ZN(_04557_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09345_ (.A1(_04468_),
    .A2(_04556_),
    .B(_04557_),
    .ZN(_01271_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09346_ (.A1(\u_cpu.rf_ram.memory[88][1] ),
    .A2(_04556_),
    .ZN(_04558_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09347_ (.A1(_04472_),
    .A2(_04556_),
    .B(_04558_),
    .ZN(_01272_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09348_ (.A1(\u_cpu.rf_ram.memory[88][2] ),
    .A2(_04556_),
    .ZN(_04559_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09349_ (.A1(_04474_),
    .A2(_04556_),
    .B(_04559_),
    .ZN(_01273_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09350_ (.A1(\u_cpu.rf_ram.memory[88][3] ),
    .A2(_04556_),
    .ZN(_04560_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09351_ (.A1(_04476_),
    .A2(_04556_),
    .B(_04560_),
    .ZN(_01274_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09352_ (.A1(\u_cpu.rf_ram.memory[88][4] ),
    .A2(_04556_),
    .ZN(_04561_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09353_ (.A1(_04478_),
    .A2(_04556_),
    .B(_04561_),
    .ZN(_01275_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09354_ (.A1(\u_cpu.rf_ram.memory[88][5] ),
    .A2(_04556_),
    .ZN(_04562_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09355_ (.A1(_04480_),
    .A2(_04556_),
    .B(_04562_),
    .ZN(_01276_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09356_ (.A1(\u_cpu.rf_ram.memory[88][6] ),
    .A2(_04556_),
    .ZN(_04563_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09357_ (.A1(_04482_),
    .A2(_04556_),
    .B(_04563_),
    .ZN(_01277_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09358_ (.A1(\u_cpu.rf_ram.memory[88][7] ),
    .A2(_04556_),
    .ZN(_04564_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09359_ (.A1(_04484_),
    .A2(_04556_),
    .B(_04564_),
    .ZN(_01278_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09360_ (.A1(_02311_),
    .A2(_01386_),
    .ZN(_04565_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09361_ (.A1(_02305_),
    .A2(_02344_),
    .A3(_02338_),
    .ZN(_04566_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09362_ (.A1(_04565_),
    .A2(_04566_),
    .Z(_04567_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09363_ (.I(_04567_),
    .Z(_04568_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09364_ (.A1(\u_cpu.cpu.genblk3.csr.o_new_irq ),
    .A2(_01392_),
    .ZN(_04569_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09365_ (.A1(_01385_),
    .A2(\u_cpu.cpu.genblk3.csr.mcause3_0[1] ),
    .ZN(_04570_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09366_ (.A1(_04569_),
    .A2(_04570_),
    .ZN(_04571_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09367_ (.A1(_04568_),
    .A2(_04571_),
    .ZN(_04572_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09368_ (.A1(_02341_),
    .A2(_04568_),
    .B(_04572_),
    .ZN(_01279_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09369_ (.A1(_01375_),
    .A2(_02306_),
    .B1(\u_cpu.cpu.genblk3.csr.mcause3_0[2] ),
    .B2(_01385_),
    .ZN(_04573_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09370_ (.A1(_04569_),
    .A2(_04573_),
    .ZN(_04574_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09371_ (.I0(_04574_),
    .I1(\u_cpu.cpu.genblk3.csr.mcause3_0[1] ),
    .S(_04568_),
    .Z(_04575_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09372_ (.I(_04575_),
    .Z(_01280_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09373_ (.A1(\u_cpu.cpu.genblk3.csr.mcause3_0[3] ),
    .A2(_01393_),
    .B(\u_cpu.cpu.genblk3.csr.o_new_irq ),
    .C(_01375_),
    .ZN(_04576_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09374_ (.A1(\u_cpu.cpu.genblk3.csr.mcause3_0[2] ),
    .A2(_04568_),
    .ZN(_04577_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09375_ (.A1(_04568_),
    .A2(_04576_),
    .B(_04577_),
    .ZN(_01281_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09376_ (.I(\u_cpu.cpu.genblk3.csr.mcause3_0[3] ),
    .ZN(_04578_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09377_ (.A1(_01381_),
    .A2(_01392_),
    .B(_04568_),
    .ZN(_04579_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09378_ (.A1(_04578_),
    .A2(_04568_),
    .B1(_04579_),
    .B2(_02349_),
    .ZN(_01282_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09379_ (.I(\u_cpu.cpu.genblk3.csr.mcause31 ),
    .ZN(_04580_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09380_ (.A1(_02311_),
    .A2(_02344_),
    .B(_01386_),
    .ZN(_04581_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09381_ (.A1(\u_cpu.cpu.genblk3.csr.o_new_irq ),
    .A2(_04581_),
    .ZN(_04582_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09382_ (.A1(_04580_),
    .A2(_04581_),
    .B1(_04582_),
    .B2(_02349_),
    .ZN(_01283_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09383_ (.I0(\u_cpu.cpu.genblk3.csr.mstatus_mie ),
    .I1(\u_cpu.cpu.genblk3.csr.mstatus_mpie ),
    .S(_04565_),
    .Z(_04583_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09384_ (.I(_04583_),
    .Z(_01284_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09385_ (.I(\u_cpu.cpu.genblk3.csr.mie_mtie ),
    .ZN(_04584_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _09386_ (.A1(\u_cpu.cpu.decode.co_ebreak ),
    .A2(\u_cpu.cpu.mem_bytecnt[1] ),
    .A3(\u_cpu.cpu.mem_bytecnt[0] ),
    .A4(_02337_),
    .ZN(_04585_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09387_ (.A1(_02339_),
    .A2(_03454_),
    .A3(_04585_),
    .ZN(_04586_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09388_ (.A1(_02348_),
    .A2(_04586_),
    .B(_01429_),
    .ZN(_04587_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09389_ (.A1(_04584_),
    .A2(_04586_),
    .B(_04587_),
    .ZN(_01285_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09390_ (.A1(_04191_),
    .A2(_02348_),
    .ZN(_04588_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09391_ (.A1(\u_cpu.cpu.genblk3.csr.mstatus_mpie ),
    .A2(_01377_),
    .B(_01393_),
    .ZN(_04589_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09392_ (.A1(_04191_),
    .A2(_02340_),
    .ZN(_04590_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09393_ (.A1(\u_cpu.cpu.genblk3.csr.mstatus_mie ),
    .A2(_04565_),
    .A3(_04590_),
    .ZN(_04591_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _09394_ (.A1(_04588_),
    .A2(_04589_),
    .A3(_04590_),
    .B(_04591_),
    .ZN(_01286_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09395_ (.A1(\u_cpu.cpu.ctrl.i_iscomp ),
    .A2(_03798_),
    .ZN(_04592_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09396_ (.A1(_03812_),
    .A2(_04592_),
    .ZN(_01287_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09397_ (.A1(\u_cpu.cpu.genblk3.csr.o_new_irq ),
    .A2(_03458_),
    .ZN(_04593_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _09398_ (.A1(_01428_),
    .A2(\u_cpu.cpu.genblk3.csr.timer_irq_r ),
    .A3(_04082_),
    .B(_04593_),
    .ZN(_01288_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09399_ (.A1(_02528_),
    .A2(_02706_),
    .ZN(_04594_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09400_ (.I(_04594_),
    .Z(_04595_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09401_ (.A1(\u_cpu.rf_ram.memory[27][0] ),
    .A2(_04595_),
    .ZN(_04596_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09402_ (.A1(_04468_),
    .A2(_04595_),
    .B(_04596_),
    .ZN(_01289_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09403_ (.A1(\u_cpu.rf_ram.memory[27][1] ),
    .A2(_04595_),
    .ZN(_04597_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09404_ (.A1(_04472_),
    .A2(_04595_),
    .B(_04597_),
    .ZN(_01290_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09405_ (.A1(\u_cpu.rf_ram.memory[27][2] ),
    .A2(_04595_),
    .ZN(_04598_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09406_ (.A1(_04474_),
    .A2(_04595_),
    .B(_04598_),
    .ZN(_01291_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09407_ (.A1(\u_cpu.rf_ram.memory[27][3] ),
    .A2(_04595_),
    .ZN(_04599_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09408_ (.A1(_04476_),
    .A2(_04595_),
    .B(_04599_),
    .ZN(_01292_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09409_ (.A1(\u_cpu.rf_ram.memory[27][4] ),
    .A2(_04595_),
    .ZN(_04600_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09410_ (.A1(_04478_),
    .A2(_04595_),
    .B(_04600_),
    .ZN(_01293_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09411_ (.A1(\u_cpu.rf_ram.memory[27][5] ),
    .A2(_04595_),
    .ZN(_04601_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09412_ (.A1(_04480_),
    .A2(_04595_),
    .B(_04601_),
    .ZN(_01294_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09413_ (.A1(\u_cpu.rf_ram.memory[27][6] ),
    .A2(_04595_),
    .ZN(_04602_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09414_ (.A1(_04482_),
    .A2(_04595_),
    .B(_04602_),
    .ZN(_01295_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09415_ (.A1(\u_cpu.rf_ram.memory[27][7] ),
    .A2(_04595_),
    .ZN(_04603_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09416_ (.A1(_04484_),
    .A2(_04595_),
    .B(_04603_),
    .ZN(_01296_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09417_ (.A1(_02528_),
    .A2(_02638_),
    .ZN(_04604_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09418_ (.I(_04604_),
    .Z(_04605_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09419_ (.A1(\u_cpu.rf_ram.memory[26][0] ),
    .A2(_04605_),
    .ZN(_04606_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09420_ (.A1(_04468_),
    .A2(_04605_),
    .B(_04606_),
    .ZN(_01297_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09421_ (.A1(\u_cpu.rf_ram.memory[26][1] ),
    .A2(_04605_),
    .ZN(_04607_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09422_ (.A1(_04472_),
    .A2(_04605_),
    .B(_04607_),
    .ZN(_01298_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09423_ (.A1(\u_cpu.rf_ram.memory[26][2] ),
    .A2(_04605_),
    .ZN(_04608_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09424_ (.A1(_04474_),
    .A2(_04605_),
    .B(_04608_),
    .ZN(_01299_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09425_ (.A1(\u_cpu.rf_ram.memory[26][3] ),
    .A2(_04605_),
    .ZN(_04609_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09426_ (.A1(_04476_),
    .A2(_04605_),
    .B(_04609_),
    .ZN(_01300_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09427_ (.A1(\u_cpu.rf_ram.memory[26][4] ),
    .A2(_04605_),
    .ZN(_04610_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09428_ (.A1(_04478_),
    .A2(_04605_),
    .B(_04610_),
    .ZN(_01301_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09429_ (.A1(\u_cpu.rf_ram.memory[26][5] ),
    .A2(_04605_),
    .ZN(_04611_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09430_ (.A1(_04480_),
    .A2(_04605_),
    .B(_04611_),
    .ZN(_01302_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09431_ (.A1(\u_cpu.rf_ram.memory[26][6] ),
    .A2(_04605_),
    .ZN(_04612_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09432_ (.A1(_04482_),
    .A2(_04605_),
    .B(_04612_),
    .ZN(_01303_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09433_ (.A1(\u_cpu.rf_ram.memory[26][7] ),
    .A2(_04605_),
    .ZN(_04613_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09434_ (.A1(_04484_),
    .A2(_04605_),
    .B(_04613_),
    .ZN(_01304_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09435_ (.A1(_02528_),
    .A2(_02695_),
    .ZN(_04614_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09436_ (.I(_04614_),
    .Z(_04615_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09437_ (.A1(\u_cpu.rf_ram.memory[25][0] ),
    .A2(_04615_),
    .ZN(_04616_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09438_ (.A1(_04468_),
    .A2(_04615_),
    .B(_04616_),
    .ZN(_01305_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09439_ (.A1(\u_cpu.rf_ram.memory[25][1] ),
    .A2(_04615_),
    .ZN(_04617_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09440_ (.A1(_04472_),
    .A2(_04615_),
    .B(_04617_),
    .ZN(_01306_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09441_ (.A1(\u_cpu.rf_ram.memory[25][2] ),
    .A2(_04615_),
    .ZN(_04618_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09442_ (.A1(_04474_),
    .A2(_04615_),
    .B(_04618_),
    .ZN(_01307_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09443_ (.A1(\u_cpu.rf_ram.memory[25][3] ),
    .A2(_04615_),
    .ZN(_04619_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09444_ (.A1(_04476_),
    .A2(_04615_),
    .B(_04619_),
    .ZN(_01308_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09445_ (.A1(\u_cpu.rf_ram.memory[25][4] ),
    .A2(_04615_),
    .ZN(_04620_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09446_ (.A1(_04478_),
    .A2(_04615_),
    .B(_04620_),
    .ZN(_01309_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09447_ (.A1(\u_cpu.rf_ram.memory[25][5] ),
    .A2(_04615_),
    .ZN(_04621_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09448_ (.A1(_04480_),
    .A2(_04615_),
    .B(_04621_),
    .ZN(_01310_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09449_ (.A1(\u_cpu.rf_ram.memory[25][6] ),
    .A2(_04615_),
    .ZN(_04622_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09450_ (.A1(_04482_),
    .A2(_04615_),
    .B(_04622_),
    .ZN(_01311_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09451_ (.A1(\u_cpu.rf_ram.memory[25][7] ),
    .A2(_04615_),
    .ZN(_04623_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09452_ (.A1(_04484_),
    .A2(_04615_),
    .B(_04623_),
    .ZN(_01312_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09453_ (.A1(_02528_),
    .A2(_02810_),
    .ZN(_04624_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09454_ (.I(_04624_),
    .Z(_04625_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09455_ (.A1(\u_cpu.rf_ram.memory[24][0] ),
    .A2(_04625_),
    .ZN(_04626_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09456_ (.A1(_04468_),
    .A2(_04625_),
    .B(_04626_),
    .ZN(_01313_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09457_ (.A1(\u_cpu.rf_ram.memory[24][1] ),
    .A2(_04625_),
    .ZN(_04627_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09458_ (.A1(_04472_),
    .A2(_04625_),
    .B(_04627_),
    .ZN(_01314_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09459_ (.A1(\u_cpu.rf_ram.memory[24][2] ),
    .A2(_04625_),
    .ZN(_04628_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09460_ (.A1(_04474_),
    .A2(_04625_),
    .B(_04628_),
    .ZN(_01315_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09461_ (.A1(\u_cpu.rf_ram.memory[24][3] ),
    .A2(_04625_),
    .ZN(_04629_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09462_ (.A1(_04476_),
    .A2(_04625_),
    .B(_04629_),
    .ZN(_01316_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09463_ (.A1(\u_cpu.rf_ram.memory[24][4] ),
    .A2(_04625_),
    .ZN(_04630_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09464_ (.A1(_04478_),
    .A2(_04625_),
    .B(_04630_),
    .ZN(_01317_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09465_ (.A1(\u_cpu.rf_ram.memory[24][5] ),
    .A2(_04625_),
    .ZN(_04631_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09466_ (.A1(_04480_),
    .A2(_04625_),
    .B(_04631_),
    .ZN(_01318_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09467_ (.A1(\u_cpu.rf_ram.memory[24][6] ),
    .A2(_04625_),
    .ZN(_04632_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09468_ (.A1(_04482_),
    .A2(_04625_),
    .B(_04632_),
    .ZN(_01319_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09469_ (.A1(\u_cpu.rf_ram.memory[24][7] ),
    .A2(_04625_),
    .ZN(_04633_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09470_ (.A1(_04484_),
    .A2(_04625_),
    .B(_04633_),
    .ZN(_01320_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09471_ (.A1(_02577_),
    .A2(_02612_),
    .ZN(_04634_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09472_ (.I0(_02573_),
    .I1(\u_cpu.rf_ram.memory[0][0] ),
    .S(_04634_),
    .Z(_04635_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09473_ (.I(_04635_),
    .Z(_01321_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09474_ (.I0(_02581_),
    .I1(\u_cpu.rf_ram.memory[0][1] ),
    .S(_04634_),
    .Z(_04636_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09475_ (.I(_04636_),
    .Z(_01322_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09476_ (.I0(_02584_),
    .I1(\u_cpu.rf_ram.memory[0][2] ),
    .S(_04634_),
    .Z(_04637_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09477_ (.I(_04637_),
    .Z(_01323_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09478_ (.I0(_02587_),
    .I1(\u_cpu.rf_ram.memory[0][3] ),
    .S(_04634_),
    .Z(_04638_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09479_ (.I(_04638_),
    .Z(_01324_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09480_ (.I0(_02590_),
    .I1(\u_cpu.rf_ram.memory[0][4] ),
    .S(_04634_),
    .Z(_04639_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09481_ (.I(_04639_),
    .Z(_01325_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09482_ (.I0(_02593_),
    .I1(\u_cpu.rf_ram.memory[0][5] ),
    .S(_04634_),
    .Z(_04640_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09483_ (.I(_04640_),
    .Z(_01326_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09484_ (.I0(_02596_),
    .I1(\u_cpu.rf_ram.memory[0][6] ),
    .S(_04634_),
    .Z(_04641_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09485_ (.I(_04641_),
    .Z(_01327_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09486_ (.I0(_02599_),
    .I1(\u_cpu.rf_ram.memory[0][7] ),
    .S(_04634_),
    .Z(_04642_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09487_ (.I(_04642_),
    .Z(_01328_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09488_ (.A1(_02469_),
    .A2(_04197_),
    .ZN(_04643_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09489_ (.I(_04643_),
    .Z(_04644_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09490_ (.A1(\u_cpu.rf_ram.memory[98][0] ),
    .A2(_04644_),
    .ZN(_04645_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09491_ (.A1(_04468_),
    .A2(_04644_),
    .B(_04645_),
    .ZN(_01329_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09492_ (.A1(\u_cpu.rf_ram.memory[98][1] ),
    .A2(_04644_),
    .ZN(_04646_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09493_ (.A1(_04472_),
    .A2(_04644_),
    .B(_04646_),
    .ZN(_01330_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09494_ (.A1(\u_cpu.rf_ram.memory[98][2] ),
    .A2(_04644_),
    .ZN(_04647_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09495_ (.A1(_04474_),
    .A2(_04644_),
    .B(_04647_),
    .ZN(_01331_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09496_ (.A1(\u_cpu.rf_ram.memory[98][3] ),
    .A2(_04644_),
    .ZN(_04648_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09497_ (.A1(_04476_),
    .A2(_04644_),
    .B(_04648_),
    .ZN(_01332_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09498_ (.A1(\u_cpu.rf_ram.memory[98][4] ),
    .A2(_04644_),
    .ZN(_04649_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09499_ (.A1(_04478_),
    .A2(_04644_),
    .B(_04649_),
    .ZN(_01333_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09500_ (.A1(\u_cpu.rf_ram.memory[98][5] ),
    .A2(_04644_),
    .ZN(_04650_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09501_ (.A1(_04480_),
    .A2(_04644_),
    .B(_04650_),
    .ZN(_01334_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09502_ (.A1(\u_cpu.rf_ram.memory[98][6] ),
    .A2(_04644_),
    .ZN(_04651_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09503_ (.A1(_04482_),
    .A2(_04644_),
    .B(_04651_),
    .ZN(_01335_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09504_ (.A1(\u_cpu.rf_ram.memory[98][7] ),
    .A2(_04644_),
    .ZN(_04652_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09505_ (.A1(_04484_),
    .A2(_04644_),
    .B(_04652_),
    .ZN(_01336_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09506_ (.A1(_02561_),
    .A2(_04197_),
    .ZN(_04653_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09507_ (.I(_04653_),
    .Z(_04654_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09508_ (.A1(\u_cpu.rf_ram.memory[100][0] ),
    .A2(_04654_),
    .ZN(_04655_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09509_ (.A1(_04468_),
    .A2(_04654_),
    .B(_04655_),
    .ZN(_01337_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09510_ (.A1(\u_cpu.rf_ram.memory[100][1] ),
    .A2(_04654_),
    .ZN(_04656_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09511_ (.A1(_04472_),
    .A2(_04654_),
    .B(_04656_),
    .ZN(_01338_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09512_ (.A1(\u_cpu.rf_ram.memory[100][2] ),
    .A2(_04654_),
    .ZN(_04657_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09513_ (.A1(_04474_),
    .A2(_04654_),
    .B(_04657_),
    .ZN(_01339_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09514_ (.A1(\u_cpu.rf_ram.memory[100][3] ),
    .A2(_04654_),
    .ZN(_04658_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09515_ (.A1(_04476_),
    .A2(_04654_),
    .B(_04658_),
    .ZN(_01340_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09516_ (.A1(\u_cpu.rf_ram.memory[100][4] ),
    .A2(_04654_),
    .ZN(_04659_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09517_ (.A1(_04478_),
    .A2(_04654_),
    .B(_04659_),
    .ZN(_01341_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09518_ (.A1(\u_cpu.rf_ram.memory[100][5] ),
    .A2(_04654_),
    .ZN(_04660_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09519_ (.A1(_04480_),
    .A2(_04654_),
    .B(_04660_),
    .ZN(_01342_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09520_ (.A1(\u_cpu.rf_ram.memory[100][6] ),
    .A2(_04654_),
    .ZN(_04661_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09521_ (.A1(_04482_),
    .A2(_04654_),
    .B(_04661_),
    .ZN(_01343_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09522_ (.A1(\u_cpu.rf_ram.memory[100][7] ),
    .A2(_04654_),
    .ZN(_04662_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09523_ (.A1(_04484_),
    .A2(_04654_),
    .B(_04662_),
    .ZN(_01344_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09524_ (.A1(_02475_),
    .A2(_02695_),
    .ZN(_04663_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09525_ (.I(_04663_),
    .Z(_04664_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09526_ (.A1(\u_cpu.rf_ram.memory[89][0] ),
    .A2(_04664_),
    .ZN(_04665_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09527_ (.A1(_04468_),
    .A2(_04664_),
    .B(_04665_),
    .ZN(_01345_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09528_ (.A1(\u_cpu.rf_ram.memory[89][1] ),
    .A2(_04664_),
    .ZN(_04666_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09529_ (.A1(_04472_),
    .A2(_04664_),
    .B(_04666_),
    .ZN(_01346_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09530_ (.A1(\u_cpu.rf_ram.memory[89][2] ),
    .A2(_04664_),
    .ZN(_04667_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09531_ (.A1(_04474_),
    .A2(_04664_),
    .B(_04667_),
    .ZN(_01347_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09532_ (.A1(\u_cpu.rf_ram.memory[89][3] ),
    .A2(_04664_),
    .ZN(_04668_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09533_ (.A1(_04476_),
    .A2(_04664_),
    .B(_04668_),
    .ZN(_01348_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09534_ (.A1(\u_cpu.rf_ram.memory[89][4] ),
    .A2(_04664_),
    .ZN(_04669_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09535_ (.A1(_04478_),
    .A2(_04664_),
    .B(_04669_),
    .ZN(_01349_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09536_ (.A1(\u_cpu.rf_ram.memory[89][5] ),
    .A2(_04664_),
    .ZN(_04670_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09537_ (.A1(_04480_),
    .A2(_04664_),
    .B(_04670_),
    .ZN(_01350_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09538_ (.A1(\u_cpu.rf_ram.memory[89][6] ),
    .A2(_04664_),
    .ZN(_04671_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09539_ (.A1(_04482_),
    .A2(_04664_),
    .B(_04671_),
    .ZN(_01351_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09540_ (.A1(\u_cpu.rf_ram.memory[89][7] ),
    .A2(_04664_),
    .ZN(_04672_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09541_ (.A1(_04484_),
    .A2(_04664_),
    .B(_04672_),
    .ZN(_01352_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09542_ (.A1(_02528_),
    .A2(_02602_),
    .ZN(_04673_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09543_ (.I(_04673_),
    .Z(_04674_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09544_ (.A1(\u_cpu.rf_ram.memory[23][0] ),
    .A2(_04674_),
    .ZN(_04675_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09545_ (.A1(_04468_),
    .A2(_04674_),
    .B(_04675_),
    .ZN(_01353_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09546_ (.A1(\u_cpu.rf_ram.memory[23][1] ),
    .A2(_04674_),
    .ZN(_04676_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09547_ (.A1(_04472_),
    .A2(_04674_),
    .B(_04676_),
    .ZN(_01354_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09548_ (.A1(\u_cpu.rf_ram.memory[23][2] ),
    .A2(_04674_),
    .ZN(_04677_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09549_ (.A1(_04474_),
    .A2(_04674_),
    .B(_04677_),
    .ZN(_01355_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09550_ (.A1(\u_cpu.rf_ram.memory[23][3] ),
    .A2(_04674_),
    .ZN(_04678_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09551_ (.A1(_04476_),
    .A2(_04674_),
    .B(_04678_),
    .ZN(_01356_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09552_ (.A1(\u_cpu.rf_ram.memory[23][4] ),
    .A2(_04674_),
    .ZN(_04679_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09553_ (.A1(_04478_),
    .A2(_04674_),
    .B(_04679_),
    .ZN(_01357_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09554_ (.A1(\u_cpu.rf_ram.memory[23][5] ),
    .A2(_04674_),
    .ZN(_04680_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09555_ (.A1(_04480_),
    .A2(_04674_),
    .B(_04680_),
    .ZN(_01358_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09556_ (.A1(\u_cpu.rf_ram.memory[23][6] ),
    .A2(_04674_),
    .ZN(_04681_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09557_ (.A1(_04482_),
    .A2(_04674_),
    .B(_04681_),
    .ZN(_01359_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09558_ (.A1(\u_cpu.rf_ram.memory[23][7] ),
    .A2(_04674_),
    .ZN(_04682_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09559_ (.A1(_04484_),
    .A2(_04674_),
    .B(_04682_),
    .ZN(_01360_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09560_ (.A1(_03797_),
    .A2(_03458_),
    .ZN(_04683_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09561_ (.A1(\u_cpu.cpu.state.ibus_cyc ),
    .A2(_04683_),
    .ZN(_04684_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09562_ (.A1(_04155_),
    .A2(_04683_),
    .B(_04684_),
    .ZN(_01361_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _09563_ (.A1(_02321_),
    .A2(_02320_),
    .A3(\u_cpu.rf_ram.rdata[7] ),
    .Z(_04685_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09564_ (.I(_04685_),
    .Z(_01362_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _09565_ (.A1(_02321_),
    .A2(\u_cpu.rf_ram.rdata[7] ),
    .A3(\u_cpu.rf_ram_if.rtrig0 ),
    .Z(_04686_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09566_ (.I(_04686_),
    .Z(_01363_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09567_ (.A1(_01429_),
    .A2(\u_cpu.rf_ram_if.rreq_r ),
    .Z(_04687_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09568_ (.I(_04687_),
    .Z(_01364_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09569_ (.A1(\u_cpu.rf_ram_if.rcnt[1] ),
    .A2(\u_cpu.rf_ram_if.rcnt[0] ),
    .Z(_04688_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09570_ (.A1(_02769_),
    .A2(_04688_),
    .ZN(_04689_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09571_ (.A1(_02783_),
    .A2(_04689_),
    .ZN(_01365_));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09572_ (.D(_00026_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[82][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09573_ (.D(_00027_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[82][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09574_ (.D(_00028_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[82][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09575_ (.D(_00029_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[82][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09576_ (.D(_00030_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[82][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09577_ (.D(_00031_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[82][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09578_ (.D(_00032_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[82][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09579_ (.D(_00033_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[82][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09580_ (.D(_00034_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[21][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09581_ (.D(_00035_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[21][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09582_ (.D(_00036_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[21][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09583_ (.D(_00037_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[21][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09584_ (.D(_00038_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[21][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09585_ (.D(_00039_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[21][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09586_ (.D(_00040_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[21][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09587_ (.D(_00041_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[21][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09588_ (.D(_00042_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[81][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09589_ (.D(_00043_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[81][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09590_ (.D(_00044_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[81][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09591_ (.D(_00045_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[81][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09592_ (.D(_00046_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[81][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09593_ (.D(_00047_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[81][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09594_ (.D(_00048_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[81][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09595_ (.D(_00049_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[81][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09596_ (.D(_00050_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[18][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09597_ (.D(_00051_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[18][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09598_ (.D(_00052_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[18][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09599_ (.D(_00053_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[18][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09600_ (.D(_00054_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[18][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09601_ (.D(_00055_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[18][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09602_ (.D(_00056_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[18][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09603_ (.D(_00057_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[18][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09604_ (.D(_00058_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[20][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09605_ (.D(_00059_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[20][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09606_ (.D(_00060_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[20][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09607_ (.D(_00061_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[20][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09608_ (.D(_00062_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[20][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09609_ (.D(_00063_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[20][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09610_ (.D(_00064_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[20][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09611_ (.D(_00065_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[20][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09612_ (.D(_00066_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[1][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09613_ (.D(_00067_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[1][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09614_ (.D(_00068_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[1][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09615_ (.D(_00069_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[1][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09616_ (.D(_00070_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[1][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09617_ (.D(_00071_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[1][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09618_ (.D(_00072_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[1][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09619_ (.D(_00073_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[1][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09620_ (.D(_00074_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[7][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09621_ (.D(_00075_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[7][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09622_ (.D(_00076_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[7][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09623_ (.D(_00077_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[7][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09624_ (.D(_00078_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[7][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09625_ (.D(_00079_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[7][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09626_ (.D(_00080_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[7][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09627_ (.D(_00081_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[7][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09628_ (.D(_00082_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[80][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09629_ (.D(_00083_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[80][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09630_ (.D(_00084_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[80][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09631_ (.D(_00085_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[80][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09632_ (.D(_00086_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[80][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09633_ (.D(_00087_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[80][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09634_ (.D(_00088_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[80][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09635_ (.D(_00089_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[80][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09636_ (.D(_00090_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[78][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09637_ (.D(_00091_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[78][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09638_ (.D(_00092_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[78][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09639_ (.D(_00093_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[78][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09640_ (.D(_00094_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[78][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09641_ (.D(_00095_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[78][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09642_ (.D(_00096_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[78][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09643_ (.D(_00097_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[78][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09644_ (.D(_00098_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[42][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09645_ (.D(_00099_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[42][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09646_ (.D(_00100_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[42][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09647_ (.D(_00101_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[42][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09648_ (.D(_00102_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[42][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09649_ (.D(_00103_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[42][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09650_ (.D(_00104_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[42][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09651_ (.D(_00105_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[42][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09652_ (.D(_00106_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[46][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09653_ (.D(_00107_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[46][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09654_ (.D(_00108_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[46][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09655_ (.D(_00109_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[46][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09656_ (.D(_00110_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[46][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09657_ (.D(_00111_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[46][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09658_ (.D(_00112_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[46][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09659_ (.D(_00113_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[46][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09660_ (.D(_00114_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[45][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09661_ (.D(_00115_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[45][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09662_ (.D(_00116_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[45][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09663_ (.D(_00117_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[45][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09664_ (.D(_00118_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[45][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09665_ (.D(_00119_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[45][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09666_ (.D(_00120_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[45][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09667_ (.D(_00121_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[45][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09668_ (.D(_00122_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[44][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09669_ (.D(_00123_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[44][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09670_ (.D(_00124_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[44][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09671_ (.D(_00125_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[44][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09672_ (.D(_00126_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[44][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09673_ (.D(_00127_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[44][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09674_ (.D(_00128_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[44][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09675_ (.D(_00129_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[44][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09676_ (.D(_00130_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[51][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09677_ (.D(_00131_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[51][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09678_ (.D(_00132_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[51][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09679_ (.D(_00133_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[51][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09680_ (.D(_00134_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[51][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09681_ (.D(_00135_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[51][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09682_ (.D(_00136_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[51][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09683_ (.D(_00137_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[51][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09684_ (.D(_00138_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[41][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09685_ (.D(_00139_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[41][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09686_ (.D(_00140_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[41][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09687_ (.D(_00141_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[41][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09688_ (.D(_00142_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[41][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09689_ (.D(_00143_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[41][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09690_ (.D(_00144_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[41][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09691_ (.D(_00145_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[41][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09692_ (.D(_00146_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[43][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09693_ (.D(_00147_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[43][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09694_ (.D(_00148_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[43][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09695_ (.D(_00149_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[43][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09696_ (.D(_00150_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[43][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09697_ (.D(_00151_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[43][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09698_ (.D(_00152_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[43][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09699_ (.D(_00153_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[43][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09700_ (.D(_00154_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[48][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09701_ (.D(_00155_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[48][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09702_ (.D(_00156_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[48][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09703_ (.D(_00157_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[48][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09704_ (.D(_00158_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[48][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09705_ (.D(_00159_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[48][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09706_ (.D(_00160_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[48][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09707_ (.D(_00161_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[48][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09708_ (.D(_00162_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[47][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09709_ (.D(_00163_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[47][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09710_ (.D(_00164_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[47][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09711_ (.D(_00165_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[47][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09712_ (.D(_00166_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[47][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09713_ (.D(_00167_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[47][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09714_ (.D(_00168_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[47][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09715_ (.D(_00169_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[47][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09716_ (.D(_00170_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[50][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09717_ (.D(_00171_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[50][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09718_ (.D(_00172_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[50][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09719_ (.D(_00173_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[50][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09720_ (.D(_00174_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[50][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09721_ (.D(_00175_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[50][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09722_ (.D(_00176_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[50][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09723_ (.D(_00177_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[50][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09724_ (.D(_00178_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[4][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09725_ (.D(_00179_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[4][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09726_ (.D(_00180_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[4][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09727_ (.D(_00181_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[4][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09728_ (.D(_00182_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[4][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09729_ (.D(_00183_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[4][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09730_ (.D(_00184_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[4][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09731_ (.D(_00185_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[4][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09732_ (.D(_00186_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram_if.rreq_r ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09733_ (.D(_00187_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram_if.rcnt[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09734_ (.D(_00188_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram_if.rcnt[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09735_ (.D(_00189_),
    .CLK(io_in[4]),
    .Q(\u_cpu.raddr[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09736_ (.D(_00190_),
    .CLK(io_in[4]),
    .Q(\u_cpu.raddr[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09737_ (.D(_00191_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[16][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09738_ (.D(_00192_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[16][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09739_ (.D(_00193_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[16][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09740_ (.D(_00194_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[16][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09741_ (.D(_00195_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[16][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09742_ (.D(_00196_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[16][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09743_ (.D(_00197_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[16][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09744_ (.D(_00198_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[16][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09745_ (.D(_00199_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[17][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09746_ (.D(_00200_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[17][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09747_ (.D(_00201_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[17][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09748_ (.D(_00202_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[17][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09749_ (.D(_00203_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[17][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09750_ (.D(_00204_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[17][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09751_ (.D(_00205_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[17][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09752_ (.D(_00206_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[17][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09753_ (.D(_00207_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[40][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09754_ (.D(_00208_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[40][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09755_ (.D(_00209_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[40][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09756_ (.D(_00210_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[40][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09757_ (.D(_00211_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[40][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09758_ (.D(_00212_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[40][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09759_ (.D(_00213_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[40][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09760_ (.D(_00214_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[40][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09761_ (.D(_00215_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[119][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09762_ (.D(_00216_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[119][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09763_ (.D(_00217_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[119][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09764_ (.D(_00218_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[119][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09765_ (.D(_00219_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[119][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09766_ (.D(_00220_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[119][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09767_ (.D(_00221_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[119][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09768_ (.D(_00222_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[119][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09769_ (.D(_00223_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[129][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09770_ (.D(_00224_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[129][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09771_ (.D(_00225_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[129][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09772_ (.D(_00226_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[129][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09773_ (.D(_00227_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[129][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09774_ (.D(_00228_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[129][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09775_ (.D(_00229_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[129][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09776_ (.D(_00230_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[129][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09777_ (.D(_00231_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[139][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09778_ (.D(_00232_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[139][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09779_ (.D(_00233_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[139][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09780_ (.D(_00234_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[139][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09781_ (.D(_00235_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[139][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09782_ (.D(_00236_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[139][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09783_ (.D(_00237_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[139][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09784_ (.D(_00238_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[139][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09785_ (.D(_00239_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[77][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09786_ (.D(_00240_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[77][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09787_ (.D(_00241_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[77][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09788_ (.D(_00242_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[77][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09789_ (.D(_00243_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[77][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09790_ (.D(_00244_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[77][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09791_ (.D(_00245_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[77][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09792_ (.D(_00246_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[77][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09793_ (.D(_00247_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[74][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09794_ (.D(_00248_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[74][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09795_ (.D(_00249_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[74][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09796_ (.D(_00250_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[74][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09797_ (.D(_00251_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[74][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09798_ (.D(_00252_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[74][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09799_ (.D(_00253_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[74][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09800_ (.D(_00254_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[74][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09801_ (.D(_00255_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[76][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09802_ (.D(_00256_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[76][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09803_ (.D(_00257_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[76][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09804_ (.D(_00258_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[76][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09805_ (.D(_00259_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[76][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09806_ (.D(_00260_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[76][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09807_ (.D(_00261_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[76][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09808_ (.D(_00262_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[76][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09809_ (.D(_00263_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[75][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09810_ (.D(_00264_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[75][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09811_ (.D(_00265_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[75][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09812_ (.D(_00266_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[75][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09813_ (.D(_00267_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[75][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09814_ (.D(_00268_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[75][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09815_ (.D(_00269_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[75][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09816_ (.D(_00270_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[75][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09817_ (.D(_00271_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[6][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09818_ (.D(_00272_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[6][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09819_ (.D(_00273_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[6][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09820_ (.D(_00274_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[6][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09821_ (.D(_00275_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[6][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09822_ (.D(_00276_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[6][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09823_ (.D(_00277_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[6][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09824_ (.D(_00278_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[6][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09825_ (.D(_00279_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[68][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09826_ (.D(_00280_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[68][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09827_ (.D(_00281_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[68][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09828_ (.D(_00282_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[68][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09829_ (.D(_00283_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[68][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09830_ (.D(_00284_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[68][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09831_ (.D(_00285_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[68][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09832_ (.D(_00286_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[68][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09833_ (.D(_00287_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[67][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09834_ (.D(_00288_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[67][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09835_ (.D(_00289_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[67][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09836_ (.D(_00290_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[67][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09837_ (.D(_00291_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[67][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09838_ (.D(_00292_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[67][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09839_ (.D(_00293_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[67][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09840_ (.D(_00294_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[67][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09841_ (.D(_00295_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[66][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09842_ (.D(_00296_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[66][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09843_ (.D(_00297_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[66][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09844_ (.D(_00298_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[66][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09845_ (.D(_00299_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[66][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09846_ (.D(_00300_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[66][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09847_ (.D(_00301_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[66][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09848_ (.D(_00302_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[66][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09849_ (.D(_00303_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[65][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09850_ (.D(_00304_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[65][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09851_ (.D(_00305_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[65][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09852_ (.D(_00306_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[65][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09853_ (.D(_00307_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[65][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09854_ (.D(_00308_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[65][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09855_ (.D(_00309_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[65][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09856_ (.D(_00310_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[65][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09857_ (.D(_00311_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[64][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09858_ (.D(_00312_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[64][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09859_ (.D(_00313_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[64][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09860_ (.D(_00314_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[64][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09861_ (.D(_00315_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[64][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09862_ (.D(_00316_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[64][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09863_ (.D(_00317_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[64][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09864_ (.D(_00318_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[64][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09865_ (.D(_00319_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[29][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09866_ (.D(_00320_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[29][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09867_ (.D(_00321_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[29][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09868_ (.D(_00322_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[29][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09869_ (.D(_00323_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[29][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09870_ (.D(_00324_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[29][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09871_ (.D(_00325_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[29][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09872_ (.D(_00326_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[29][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09873_ (.D(_00327_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[63][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09874_ (.D(_00328_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[63][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09875_ (.D(_00329_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[63][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09876_ (.D(_00330_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[63][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09877_ (.D(_00331_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[63][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09878_ (.D(_00332_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[63][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09879_ (.D(_00333_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[63][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09880_ (.D(_00334_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[63][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09881_ (.D(_00335_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[62][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09882_ (.D(_00336_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[62][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09883_ (.D(_00337_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[62][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09884_ (.D(_00338_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[62][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09885_ (.D(_00339_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[62][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09886_ (.D(_00340_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[62][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09887_ (.D(_00341_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[62][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09888_ (.D(_00342_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[62][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09889_ (.D(_00343_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[61][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09890_ (.D(_00344_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[61][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09891_ (.D(_00345_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[61][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09892_ (.D(_00346_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[61][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09893_ (.D(_00347_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[61][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09894_ (.D(_00348_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[61][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09895_ (.D(_00349_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[61][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09896_ (.D(_00350_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[61][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09897_ (.D(_00351_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[60][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09898_ (.D(_00352_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[60][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09899_ (.D(_00353_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[60][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09900_ (.D(_00354_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[60][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09901_ (.D(_00355_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[60][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09902_ (.D(_00356_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[60][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09903_ (.D(_00357_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[60][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09904_ (.D(_00358_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[60][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09905_ (.D(_00359_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[19][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09906_ (.D(_00360_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[19][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09907_ (.D(_00361_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[19][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09908_ (.D(_00362_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[19][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09909_ (.D(_00363_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[19][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09910_ (.D(_00364_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[19][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09911_ (.D(_00365_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[19][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09912_ (.D(_00366_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[19][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09913_ (.D(_00367_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[5][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09914_ (.D(_00368_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[5][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09915_ (.D(_00369_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[5][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09916_ (.D(_00370_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[5][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09917_ (.D(_00371_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[5][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09918_ (.D(_00372_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[5][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09919_ (.D(_00373_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[5][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09920_ (.D(_00374_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[5][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09921_ (.D(_00375_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[58][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09922_ (.D(_00376_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[58][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09923_ (.D(_00377_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[58][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09924_ (.D(_00378_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[58][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09925_ (.D(_00379_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[58][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09926_ (.D(_00380_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[58][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09927_ (.D(_00381_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[58][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09928_ (.D(_00382_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[58][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09929_ (.D(_00383_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[57][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09930_ (.D(_00384_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[57][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09931_ (.D(_00385_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[57][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09932_ (.D(_00386_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[57][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09933_ (.D(_00387_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[57][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09934_ (.D(_00388_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[57][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09935_ (.D(_00389_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[57][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09936_ (.D(_00390_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[57][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09937_ (.D(_00391_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[56][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09938_ (.D(_00392_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[56][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09939_ (.D(_00393_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[56][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09940_ (.D(_00394_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[56][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09941_ (.D(_00395_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[56][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09942_ (.D(_00396_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[56][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09943_ (.D(_00397_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[56][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09944_ (.D(_00398_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[56][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09945_ (.D(_00399_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[55][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09946_ (.D(_00400_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[55][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09947_ (.D(_00401_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[55][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09948_ (.D(_00402_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[55][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09949_ (.D(_00403_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[55][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09950_ (.D(_00404_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[55][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09951_ (.D(_00405_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[55][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09952_ (.D(_00406_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[55][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09953_ (.D(_00407_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[54][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09954_ (.D(_00408_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[54][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09955_ (.D(_00409_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[54][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09956_ (.D(_00410_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[54][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09957_ (.D(_00411_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[54][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09958_ (.D(_00412_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[54][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09959_ (.D(_00413_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[54][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09960_ (.D(_00414_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[54][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09961_ (.D(_00415_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[53][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09962_ (.D(_00416_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[53][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09963_ (.D(_00417_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[53][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09964_ (.D(_00418_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[53][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09965_ (.D(_00419_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[53][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09966_ (.D(_00420_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[53][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09967_ (.D(_00421_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[53][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09968_ (.D(_00422_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[53][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09969_ (.D(_00423_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[52][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09970_ (.D(_00424_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[52][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09971_ (.D(_00425_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[52][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09972_ (.D(_00426_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[52][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09973_ (.D(_00427_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[52][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09974_ (.D(_00428_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[52][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09975_ (.D(_00429_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[52][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09976_ (.D(_00430_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[52][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09977_ (.D(_00431_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[9][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09978_ (.D(_00432_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[9][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09979_ (.D(_00433_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[9][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09980_ (.D(_00434_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[9][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09981_ (.D(_00435_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[9][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09982_ (.D(_00436_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[9][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09983_ (.D(_00437_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[9][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09984_ (.D(_00438_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[9][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09985_ (.D(_00439_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[15][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09986_ (.D(_00440_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[15][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09987_ (.D(_00441_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[15][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09988_ (.D(_00442_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[15][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09989_ (.D(_00443_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[15][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09990_ (.D(_00444_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[15][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09991_ (.D(_00445_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[15][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09992_ (.D(_00446_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[15][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09993_ (.D(_00000_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.rdata[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09994_ (.D(_00001_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.rdata[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09995_ (.D(_00002_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.rdata[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09996_ (.D(_00003_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.rdata[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09997_ (.D(_00004_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.rdata[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09998_ (.D(_00005_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.rdata[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _09999_ (.D(_00006_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.rdata[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10000_ (.D(_00007_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.rdata[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10001_ (.D(_00447_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[142][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10002_ (.D(_00448_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[142][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10003_ (.D(_00449_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[142][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10004_ (.D(_00450_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[142][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10005_ (.D(_00451_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[142][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10006_ (.D(_00452_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[142][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10007_ (.D(_00453_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[142][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10008_ (.D(_00454_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[142][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10009_ (.D(_00455_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[141][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10010_ (.D(_00456_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[141][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10011_ (.D(_00457_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[141][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10012_ (.D(_00458_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[141][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10013_ (.D(_00459_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[141][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10014_ (.D(_00460_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[141][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10015_ (.D(_00461_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[141][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10016_ (.D(_00462_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[141][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10017_ (.D(_00463_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[140][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10018_ (.D(_00464_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[140][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10019_ (.D(_00465_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[140][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10020_ (.D(_00466_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[140][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10021_ (.D(_00467_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[140][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10022_ (.D(_00468_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[140][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10023_ (.D(_00469_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[140][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10024_ (.D(_00470_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[140][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10025_ (.D(_00471_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[13][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10026_ (.D(_00472_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[13][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10027_ (.D(_00473_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[13][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10028_ (.D(_00474_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[13][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10029_ (.D(_00475_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[13][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10030_ (.D(_00476_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[13][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10031_ (.D(_00477_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[13][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10032_ (.D(_00478_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[13][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10033_ (.D(_00479_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[72][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10034_ (.D(_00480_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[72][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10035_ (.D(_00481_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[72][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10036_ (.D(_00482_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[72][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10037_ (.D(_00483_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[72][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10038_ (.D(_00484_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[72][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10039_ (.D(_00485_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[72][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10040_ (.D(_00486_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[72][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10041_ (.D(_00487_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[73][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10042_ (.D(_00488_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[73][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10043_ (.D(_00489_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[73][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10044_ (.D(_00490_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[73][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10045_ (.D(_00491_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[73][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10046_ (.D(_00492_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[73][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10047_ (.D(_00493_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[73][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10048_ (.D(_00494_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[73][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10049_ (.D(_00495_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[71][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10050_ (.D(_00496_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[71][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10051_ (.D(_00497_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[71][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10052_ (.D(_00498_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[71][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10053_ (.D(_00499_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[71][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10054_ (.D(_00500_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[71][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10055_ (.D(_00501_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[71][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10056_ (.D(_00502_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[71][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10057_ (.D(_00503_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[70][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10058_ (.D(_00504_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[70][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10059_ (.D(_00505_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[70][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10060_ (.D(_00506_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[70][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10061_ (.D(_00507_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[70][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10062_ (.D(_00508_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[70][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10063_ (.D(_00509_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[70][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10064_ (.D(_00510_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[70][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10065_ (.D(_00511_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[143][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10066_ (.D(_00512_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[143][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10067_ (.D(_00513_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[143][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10068_ (.D(_00514_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[143][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10069_ (.D(_00515_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[143][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10070_ (.D(_00516_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[143][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10071_ (.D(_00517_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[143][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10072_ (.D(_00518_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[143][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10073_ (.D(_00519_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[14][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10074_ (.D(_00520_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[14][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10075_ (.D(_00521_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[14][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10076_ (.D(_00522_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[14][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10077_ (.D(_00523_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[14][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10078_ (.D(_00524_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[14][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10079_ (.D(_00525_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[14][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10080_ (.D(_00526_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[14][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10081_ (.D(_00527_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[138][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10082_ (.D(_00528_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[138][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10083_ (.D(_00529_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[138][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10084_ (.D(_00530_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[138][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10085_ (.D(_00531_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[138][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10086_ (.D(_00532_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[138][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10087_ (.D(_00533_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[138][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10088_ (.D(_00534_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[138][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10089_ (.D(_00535_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[39][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10090_ (.D(_00536_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[39][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10091_ (.D(_00537_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[39][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10092_ (.D(_00538_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[39][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10093_ (.D(_00539_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[39][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10094_ (.D(_00540_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[39][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10095_ (.D(_00541_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[39][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10096_ (.D(_00542_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[39][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10097_ (.D(_00543_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[137][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10098_ (.D(_00544_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[137][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10099_ (.D(_00545_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[137][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10100_ (.D(_00546_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[137][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10101_ (.D(_00547_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[137][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10102_ (.D(_00548_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[137][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10103_ (.D(_00549_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[137][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10104_ (.D(_00550_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[137][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10105_ (.D(_00551_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[49][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10106_ (.D(_00552_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[49][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10107_ (.D(_00553_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[49][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10108_ (.D(_00554_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[49][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10109_ (.D(_00555_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[49][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10110_ (.D(_00556_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[49][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10111_ (.D(_00557_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[49][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10112_ (.D(_00558_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[49][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10113_ (.D(_00559_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[136][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10114_ (.D(_00560_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[136][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10115_ (.D(_00561_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[136][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10116_ (.D(_00562_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[136][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10117_ (.D(_00563_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[136][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10118_ (.D(_00564_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[136][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10119_ (.D(_00565_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[136][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10120_ (.D(_00566_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[136][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10121_ (.D(_00567_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[135][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10122_ (.D(_00568_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[135][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10123_ (.D(_00569_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[135][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10124_ (.D(_00570_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[135][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10125_ (.D(_00571_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[135][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10126_ (.D(_00572_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[135][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10127_ (.D(_00573_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[135][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10128_ (.D(_00574_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[135][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10129_ (.D(_00575_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[134][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10130_ (.D(_00576_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[134][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10131_ (.D(_00577_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[134][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10132_ (.D(_00578_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[134][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10133_ (.D(_00579_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[134][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10134_ (.D(_00580_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[134][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10135_ (.D(_00581_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[134][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10136_ (.D(_00582_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[134][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10137_ (.D(_00583_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[133][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10138_ (.D(_00584_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[133][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10139_ (.D(_00585_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[133][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10140_ (.D(_00586_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[133][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10141_ (.D(_00587_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[133][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10142_ (.D(_00588_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[133][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10143_ (.D(_00589_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[133][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10144_ (.D(_00590_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[133][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10145_ (.D(_00591_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[132][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10146_ (.D(_00592_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[132][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10147_ (.D(_00593_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[132][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10148_ (.D(_00594_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[132][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10149_ (.D(_00595_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[132][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10150_ (.D(_00596_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[132][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10151_ (.D(_00597_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[132][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10152_ (.D(_00598_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[132][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10153_ (.D(_00599_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[131][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10154_ (.D(_00600_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[131][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10155_ (.D(_00601_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[131][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10156_ (.D(_00602_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[131][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10157_ (.D(_00603_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[131][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10158_ (.D(_00604_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[131][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10159_ (.D(_00605_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[131][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10160_ (.D(_00606_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[131][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10161_ (.D(_00607_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[130][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10162_ (.D(_00608_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[130][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10163_ (.D(_00609_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[130][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10164_ (.D(_00610_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[130][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10165_ (.D(_00611_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[130][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10166_ (.D(_00612_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[130][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10167_ (.D(_00613_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[130][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10168_ (.D(_00614_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[130][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10169_ (.D(_00615_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[12][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10170_ (.D(_00616_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[12][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10171_ (.D(_00617_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[12][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10172_ (.D(_00618_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[12][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10173_ (.D(_00619_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[12][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10174_ (.D(_00620_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[12][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10175_ (.D(_00621_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[12][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10176_ (.D(_00622_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[12][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10177_ (.D(_00623_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[22][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10178_ (.D(_00624_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[22][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10179_ (.D(_00625_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[22][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10180_ (.D(_00626_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[22][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10181_ (.D(_00627_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[22][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10182_ (.D(_00628_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[22][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10183_ (.D(_00629_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[22][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10184_ (.D(_00630_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[22][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10185_ (.D(_00631_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[128][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10186_ (.D(_00632_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[128][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10187_ (.D(_00633_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[128][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10188_ (.D(_00634_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[128][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10189_ (.D(_00635_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[128][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10190_ (.D(_00636_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[128][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10191_ (.D(_00637_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[128][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10192_ (.D(_00638_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[128][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10193_ (.D(_00639_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[127][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10194_ (.D(_00640_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[127][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10195_ (.D(_00641_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[127][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10196_ (.D(_00642_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[127][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10197_ (.D(_00643_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[127][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10198_ (.D(_00644_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[127][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10199_ (.D(_00645_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[127][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10200_ (.D(_00646_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[127][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10201_ (.D(_00647_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[126][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10202_ (.D(_00648_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[126][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10203_ (.D(_00649_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[126][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10204_ (.D(_00650_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[126][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10205_ (.D(_00651_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[126][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10206_ (.D(_00652_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[126][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10207_ (.D(_00653_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[126][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10208_ (.D(_00654_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[126][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10209_ (.D(_00655_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[125][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10210_ (.D(_00656_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[125][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10211_ (.D(_00657_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[125][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10212_ (.D(_00658_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[125][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10213_ (.D(_00659_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[125][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10214_ (.D(_00660_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[125][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10215_ (.D(_00661_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[125][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10216_ (.D(_00662_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[125][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10217_ (.D(_00663_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[124][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10218_ (.D(_00664_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[124][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10219_ (.D(_00665_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[124][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10220_ (.D(_00666_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[124][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10221_ (.D(_00667_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[124][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10222_ (.D(_00668_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[124][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10223_ (.D(_00669_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[124][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10224_ (.D(_00670_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[124][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10225_ (.D(_00015_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram_if.rdata1[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10226_ (.D(_00016_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram_if.rdata1[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10227_ (.D(_00017_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram_if.rdata1[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10228_ (.D(_00018_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram_if.rdata1[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10229_ (.D(_00019_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram_if.rdata1[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10230_ (.D(_00020_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram_if.rdata1[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10231_ (.D(_00671_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[123][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10232_ (.D(_00672_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[123][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10233_ (.D(_00673_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[123][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10234_ (.D(_00674_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[123][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10235_ (.D(_00675_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[123][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10236_ (.D(_00676_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[123][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10237_ (.D(_00677_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[123][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10238_ (.D(_00678_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[123][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10239_ (.D(_00008_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.alu.i_rs1 ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10240_ (.D(_00009_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram_if.rdata0[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10241_ (.D(_00010_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram_if.rdata0[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10242_ (.D(_00011_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram_if.rdata0[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10243_ (.D(_00012_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram_if.rdata0[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10244_ (.D(_00013_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram_if.rdata0[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10245_ (.D(_00014_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram_if.rdata0[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10246_ (.D(_00679_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[38][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10247_ (.D(_00680_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[38][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10248_ (.D(_00681_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[38][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10249_ (.D(_00682_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[38][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10250_ (.D(_00683_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[38][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10251_ (.D(_00684_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[38][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10252_ (.D(_00685_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[38][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10253_ (.D(_00686_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[38][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10254_ (.D(_00687_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[37][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10255_ (.D(_00688_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[37][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10256_ (.D(_00689_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[37][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10257_ (.D(_00690_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[37][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10258_ (.D(_00691_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[37][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10259_ (.D(_00692_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[37][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10260_ (.D(_00693_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[37][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10261_ (.D(_00694_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[37][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10262_ (.D(_00695_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[36][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10263_ (.D(_00696_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[36][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10264_ (.D(_00697_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[36][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10265_ (.D(_00698_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[36][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10266_ (.D(_00699_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[36][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10267_ (.D(_00700_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[36][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10268_ (.D(_00701_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[36][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10269_ (.D(_00702_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[36][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10270_ (.D(_00703_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.state.stage_two_req ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10271_ (.D(_00704_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.state.o_cnt[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10272_ (.D(_00705_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.mem_bytecnt[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10273_ (.D(_00706_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.mem_bytecnt[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10274_ (.D(_00707_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.state.o_cnt_r[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10275_ (.D(_00708_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.state.o_cnt_r[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10276_ (.D(_00709_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.state.o_cnt_r[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10277_ (.D(_00710_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.state.o_cnt_r[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10278_ (.D(_00711_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[91][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10279_ (.D(_00712_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[91][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10280_ (.D(_00713_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[91][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10281_ (.D(_00714_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[91][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10282_ (.D(_00715_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[91][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10283_ (.D(_00716_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[91][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10284_ (.D(_00717_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[91][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10285_ (.D(_00718_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[91][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10286_ (.D(_00719_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[90][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10287_ (.D(_00720_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[90][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10288_ (.D(_00721_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[90][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10289_ (.D(_00722_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[90][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10290_ (.D(_00723_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[90][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10291_ (.D(_00724_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[90][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10292_ (.D(_00725_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[90][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10293_ (.D(_00726_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[90][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10294_ (.D(_00727_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.state.genblk1.misalign_trap_sync_r ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10295_ (.D(_00728_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.mem_if.signbit ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10296_ (.D(_00729_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.ctrl.i_jump ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10297_ (.D(_00730_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.bufreg2.i_cnt_done ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10298_ (.D(_00731_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.state.init_done ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10299_ (.D(_00732_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[92][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10300_ (.D(_00733_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[92][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10301_ (.D(_00734_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[92][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10302_ (.D(_00735_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[92][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10303_ (.D(_00736_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[92][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10304_ (.D(_00737_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[92][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10305_ (.D(_00738_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[92][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10306_ (.D(_00739_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[92][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10307_ (.D(_00740_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[35][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10308_ (.D(_00741_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[35][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10309_ (.D(_00742_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[35][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10310_ (.D(_00743_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[35][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10311_ (.D(_00744_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[35][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10312_ (.D(_00745_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[35][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10313_ (.D(_00746_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[35][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10314_ (.D(_00747_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[35][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10315_ (.D(_00748_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[34][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10316_ (.D(_00749_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[34][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10317_ (.D(_00750_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[34][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10318_ (.D(_00751_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[34][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10319_ (.D(_00752_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[34][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10320_ (.D(_00753_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[34][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10321_ (.D(_00754_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[34][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10322_ (.D(_00755_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[34][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10323_ (.D(_00756_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[117][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10324_ (.D(_00757_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[117][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10325_ (.D(_00758_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[117][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10326_ (.D(_00759_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[117][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10327_ (.D(_00760_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[117][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10328_ (.D(_00761_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[117][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10329_ (.D(_00762_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[117][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10330_ (.D(_00763_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[117][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10331_ (.D(_00764_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[120][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10332_ (.D(_00765_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[120][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10333_ (.D(_00766_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[120][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10334_ (.D(_00767_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[120][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10335_ (.D(_00768_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[120][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10336_ (.D(_00769_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[120][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10337_ (.D(_00770_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[120][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10338_ (.D(_00771_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[120][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10339_ (.D(_00772_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[118][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10340_ (.D(_00773_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[118][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10341_ (.D(_00774_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[118][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10342_ (.D(_00775_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[118][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10343_ (.D(_00776_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[118][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10344_ (.D(_00777_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[118][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10345_ (.D(_00778_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[118][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10346_ (.D(_00779_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[118][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10347_ (.D(_00780_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[121][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10348_ (.D(_00781_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[121][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10349_ (.D(_00782_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[121][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10350_ (.D(_00783_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[121][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10351_ (.D(_00784_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[121][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10352_ (.D(_00785_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[121][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10353_ (.D(_00786_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[121][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10354_ (.D(_00787_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[121][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10355_ (.D(_00788_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[8][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10356_ (.D(_00789_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[8][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10357_ (.D(_00790_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[8][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10358_ (.D(_00791_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[8][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10359_ (.D(_00792_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[8][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10360_ (.D(_00793_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[8][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10361_ (.D(_00794_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[8][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10362_ (.D(_00795_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[8][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10363_ (.D(_00796_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[11][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10364_ (.D(_00797_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[11][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10365_ (.D(_00798_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[11][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10366_ (.D(_00799_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[11][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10367_ (.D(_00800_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[11][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10368_ (.D(_00801_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[11][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10369_ (.D(_00802_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[11][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10370_ (.D(_00803_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[11][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10371_ (.D(_00804_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[112][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10372_ (.D(_00805_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[112][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10373_ (.D(_00806_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[112][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10374_ (.D(_00807_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[112][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10375_ (.D(_00808_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[112][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10376_ (.D(_00809_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[112][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10377_ (.D(_00810_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[112][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10378_ (.D(_00811_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[112][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10379_ (.D(_00812_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[122][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10380_ (.D(_00813_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[122][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10381_ (.D(_00814_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[122][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10382_ (.D(_00815_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[122][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10383_ (.D(_00816_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[122][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10384_ (.D(_00817_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[122][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10385_ (.D(_00818_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[122][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10386_ (.D(_00819_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[122][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10387_ (.D(_00820_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[115][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10388_ (.D(_00821_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[115][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10389_ (.D(_00822_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[115][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10390_ (.D(_00823_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[115][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10391_ (.D(_00824_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[115][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10392_ (.D(_00825_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[115][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10393_ (.D(_00826_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[115][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10394_ (.D(_00827_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[115][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10395_ (.D(_00828_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[116][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10396_ (.D(_00829_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[116][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10397_ (.D(_00830_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[116][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10398_ (.D(_00831_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[116][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10399_ (.D(_00832_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[116][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10400_ (.D(_00833_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[116][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10401_ (.D(_00834_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[116][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10402_ (.D(_00835_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[116][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10403_ (.D(_00836_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[33][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10404_ (.D(_00837_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[33][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10405_ (.D(_00838_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[33][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10406_ (.D(_00839_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[33][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10407_ (.D(_00840_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[33][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10408_ (.D(_00841_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[33][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10409_ (.D(_00842_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[33][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10410_ (.D(_00843_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[33][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10411_ (.D(_00844_),
    .CLK(io_in[4]),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10412_ (.D(_00845_),
    .CLK(io_in[4]),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10413_ (.D(_00846_),
    .CLK(io_in[4]),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10414_ (.D(_00847_),
    .CLK(io_in[4]),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10415_ (.D(_00848_),
    .CLK(io_in[4]),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10416_ (.D(_00849_),
    .CLK(io_in[4]),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10417_ (.D(_00850_),
    .CLK(io_in[4]),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10418_ (.D(_00851_),
    .CLK(io_in[4]),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10419_ (.D(_00852_),
    .CLK(io_in[4]),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10420_ (.D(_00853_),
    .CLK(io_in[4]),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10421_ (.D(_00854_),
    .CLK(io_in[4]),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10422_ (.D(_00855_),
    .CLK(io_in[4]),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10423_ (.D(_00856_),
    .CLK(io_in[4]),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10424_ (.D(_00857_),
    .CLK(io_in[4]),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10425_ (.D(_00858_),
    .CLK(io_in[4]),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10426_ (.D(_00859_),
    .CLK(io_in[4]),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10427_ (.D(_00860_),
    .CLK(io_in[4]),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10428_ (.D(_00861_),
    .CLK(io_in[4]),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10429_ (.D(_00862_),
    .CLK(io_in[4]),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10430_ (.D(_00863_),
    .CLK(io_in[4]),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10431_ (.D(_00864_),
    .CLK(io_in[4]),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10432_ (.D(_00865_),
    .CLK(io_in[4]),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10433_ (.D(_00866_),
    .CLK(io_in[4]),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10434_ (.D(_00867_),
    .CLK(io_in[4]),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10435_ (.D(_00868_),
    .CLK(io_in[4]),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10436_ (.D(_00869_),
    .CLK(io_in[4]),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10437_ (.D(_00870_),
    .CLK(io_in[4]),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10438_ (.D(_00871_),
    .CLK(io_in[4]),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10439_ (.D(_00872_),
    .CLK(io_in[4]),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10440_ (.D(_00873_),
    .CLK(io_in[4]),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[29] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10441_ (.D(_00874_),
    .CLK(io_in[4]),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[30] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10442_ (.D(_00875_),
    .CLK(io_in[4]),
    .Q(\u_arbiter.i_wb_cpu_dbus_dat[31] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10443_ (.D(_00876_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[113][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10444_ (.D(_00877_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[113][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10445_ (.D(_00878_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[113][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10446_ (.D(_00879_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[113][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10447_ (.D(_00880_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[113][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10448_ (.D(_00881_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[113][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10449_ (.D(_00882_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[113][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10450_ (.D(_00883_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[113][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10451_ (.D(_00884_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.decode.opcode[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10452_ (.D(_00885_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.decode.opcode[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10453_ (.D(_00886_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.decode.opcode[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10454_ (.D(_00887_),
    .CLK(io_in[4]),
    .Q(\u_arbiter.i_wb_cpu_dbus_we ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10455_ (.D(_00888_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.branch_op ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10456_ (.D(_00889_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.bne_or_bge ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10457_ (.D(_00890_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.decode.co_mem_word ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10458_ (.D(_00891_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.csr_d_sel ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10459_ (.D(_00892_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.decode.co_ebreak ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10460_ (.D(_00893_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.decode.op21 ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10461_ (.D(_00894_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.decode.op22 ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10462_ (.D(_00895_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[114][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10463_ (.D(_00896_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[114][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10464_ (.D(_00897_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[114][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10465_ (.D(_00898_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[114][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10466_ (.D(_00899_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[114][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10467_ (.D(_00900_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[114][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10468_ (.D(_00901_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[114][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10469_ (.D(_00902_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[114][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10470_ (.D(_00903_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.decode.op26 ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10471_ (.D(_00904_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.immdec.imm24_20[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10472_ (.D(_00905_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.immdec.imm24_20[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10473_ (.D(_00906_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.immdec.imm24_20[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10474_ (.D(_00907_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.immdec.imm24_20[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10475_ (.D(_00908_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.immdec.imm24_20[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10476_ (.D(_00909_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.immdec.imm30_25[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10477_ (.D(_00910_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.immdec.imm30_25[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10478_ (.D(_00911_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.immdec.imm30_25[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10479_ (.D(_00912_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.immdec.imm30_25[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10480_ (.D(_00913_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.immdec.imm30_25[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10481_ (.D(_00914_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.immdec.imm30_25[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10482_ (.D(_00915_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.immdec.imm7 ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10483_ (.D(_00916_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.immdec.imm19_12_20[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10484_ (.D(_00917_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.immdec.imm19_12_20[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10485_ (.D(_00918_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.immdec.imm19_12_20[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10486_ (.D(_00919_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.immdec.imm19_12_20[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10487_ (.D(_00920_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.csr_imm ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10488_ (.D(_00921_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.immdec.imm19_12_20[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10489_ (.D(_00922_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.immdec.imm19_12_20[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10490_ (.D(_00923_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.immdec.imm19_12_20[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10491_ (.D(_00924_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.immdec.imm19_12_20[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10492_ (.D(_00925_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.immdec.imm31 ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10493_ (.D(_00926_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.genblk3.csr.timer_irq_r ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10494_ (.D(_00927_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[32][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10495_ (.D(_00928_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[32][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10496_ (.D(_00929_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[32][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10497_ (.D(_00930_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[32][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10498_ (.D(_00931_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[32][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10499_ (.D(_00932_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[32][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10500_ (.D(_00933_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[32][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10501_ (.D(_00934_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[32][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10502_ (.D(_00935_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[31][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10503_ (.D(_00936_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[31][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10504_ (.D(_00937_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[31][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10505_ (.D(_00938_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[31][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10506_ (.D(_00939_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[31][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10507_ (.D(_00940_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[31][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10508_ (.D(_00941_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[31][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10509_ (.D(_00942_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[31][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10510_ (.D(_00943_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.alu.cmp_r ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10511_ (.D(_00944_),
    .CLK(io_in[4]),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10512_ (.D(_00945_),
    .CLK(io_in[4]),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10513_ (.D(_00946_),
    .CLK(io_in[4]),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10514_ (.D(_00947_),
    .CLK(io_in[4]),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10515_ (.D(_00948_),
    .CLK(io_in[4]),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10516_ (.D(_00949_),
    .CLK(io_in[4]),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10517_ (.D(_00950_),
    .CLK(io_in[4]),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10518_ (.D(_00951_),
    .CLK(io_in[4]),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10519_ (.D(_00952_),
    .CLK(io_in[4]),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10520_ (.D(_00953_),
    .CLK(io_in[4]),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10521_ (.D(_00954_),
    .CLK(io_in[4]),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10522_ (.D(_00955_),
    .CLK(io_in[4]),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10523_ (.D(_00956_),
    .CLK(io_in[4]),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10524_ (.D(_00957_),
    .CLK(io_in[4]),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10525_ (.D(_00958_),
    .CLK(io_in[4]),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10526_ (.D(_00959_),
    .CLK(io_in[4]),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10527_ (.D(_00960_),
    .CLK(io_in[4]),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10528_ (.D(_00961_),
    .CLK(io_in[4]),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10529_ (.D(_00962_),
    .CLK(io_in[4]),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10530_ (.D(_00963_),
    .CLK(io_in[4]),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10531_ (.D(_00964_),
    .CLK(io_in[4]),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10532_ (.D(_00965_),
    .CLK(io_in[4]),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10533_ (.D(_00966_),
    .CLK(io_in[4]),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10534_ (.D(_00967_),
    .CLK(io_in[4]),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10535_ (.D(_00968_),
    .CLK(io_in[4]),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10536_ (.D(_00969_),
    .CLK(io_in[4]),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10537_ (.D(_00970_),
    .CLK(io_in[4]),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10538_ (.D(_00971_),
    .CLK(io_in[4]),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[29] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10539_ (.D(_00972_),
    .CLK(io_in[4]),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[30] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10540_ (.D(_00973_),
    .CLK(io_in[4]),
    .Q(\u_arbiter.i_wb_cpu_dbus_adr[31] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10541_ (.D(_00022_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.bufreg.c_r ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10542_ (.D(_00974_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.bufreg.lsb[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10543_ (.D(_00975_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.bufreg.lsb[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10544_ (.D(_00976_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[30][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10545_ (.D(_00977_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[30][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10546_ (.D(_00978_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[30][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10547_ (.D(_00979_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[30][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10548_ (.D(_00980_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[30][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10549_ (.D(_00981_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[30][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10550_ (.D(_00982_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[30][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10551_ (.D(_00983_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[30][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10552_ (.D(_00024_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.ctrl.pc_plus_offset_cy_r ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10553_ (.D(_00023_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.ctrl.pc_plus_4_cy_r ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10554_ (.D(_00984_),
    .CLK(io_in[4]),
    .Q(\u_arbiter.i_wb_cpu_ibus_adr[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10555_ (.D(_00985_),
    .CLK(io_in[4]),
    .Q(\u_arbiter.i_wb_cpu_ibus_adr[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10556_ (.D(_00986_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10557_ (.D(_00987_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10558_ (.D(_00988_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10559_ (.D(_00989_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10560_ (.D(_00990_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10561_ (.D(_00991_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10562_ (.D(_00992_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10563_ (.D(_00993_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10564_ (.D(_00994_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10565_ (.D(_00995_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10566_ (.D(_00996_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10567_ (.D(_00997_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10568_ (.D(_00998_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10569_ (.D(_00999_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10570_ (.D(_01000_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10571_ (.D(_01001_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10572_ (.D(_01002_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10573_ (.D(_01003_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10574_ (.D(_01004_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10575_ (.D(_01005_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10576_ (.D(_01006_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10577_ (.D(_01007_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10578_ (.D(_01008_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10579_ (.D(_01009_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10580_ (.D(_01010_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10581_ (.D(_01011_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10582_ (.D(_01012_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10583_ (.D(_01013_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[29] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10584_ (.D(_01014_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[30] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10585_ (.D(_01015_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.ctrl.o_ibus_adr[31] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10586_ (.D(_01016_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[109][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10587_ (.D(_01017_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[109][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10588_ (.D(_01018_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[109][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10589_ (.D(_01019_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[109][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10590_ (.D(_01020_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[109][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10591_ (.D(_01021_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[109][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10592_ (.D(_01022_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[109][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10593_ (.D(_01023_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[109][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10594_ (.D(_00021_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.alu.add_cy_r ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10595_ (.D(_01024_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[3][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10596_ (.D(_01025_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[3][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10597_ (.D(_01026_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[3][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10598_ (.D(_01027_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[3][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10599_ (.D(_01028_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[3][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10600_ (.D(_01029_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[3][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10601_ (.D(_01030_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[3][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10602_ (.D(_01031_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[3][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10603_ (.D(_01032_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[2][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10604_ (.D(_01033_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[2][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10605_ (.D(_01034_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[2][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10606_ (.D(_01035_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[2][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10607_ (.D(_01036_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[2][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10608_ (.D(_01037_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[2][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10609_ (.D(_01038_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[2][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10610_ (.D(_01039_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[2][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10611_ (.D(_01040_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[93][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10612_ (.D(_01041_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[93][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10613_ (.D(_01042_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[93][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10614_ (.D(_01043_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[93][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10615_ (.D(_01044_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[93][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10616_ (.D(_01045_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[93][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10617_ (.D(_01046_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[93][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10618_ (.D(_01047_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[93][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10619_ (.D(_01048_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.immdec.imm11_7[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10620_ (.D(_01049_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.immdec.imm11_7[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10621_ (.D(_01050_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.immdec.imm11_7[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10622_ (.D(_01051_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.immdec.imm11_7[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10623_ (.D(_01052_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.immdec.imm11_7[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10624_ (.D(_01053_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[97][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10625_ (.D(_01054_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[97][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10626_ (.D(_01055_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[97][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10627_ (.D(_01056_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[97][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10628_ (.D(_01057_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[97][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10629_ (.D(_01058_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[97][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10630_ (.D(_01059_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[97][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10631_ (.D(_01060_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[97][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10632_ (.D(_01061_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[94][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10633_ (.D(_01062_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[94][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10634_ (.D(_01063_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[94][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10635_ (.D(_01064_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[94][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10636_ (.D(_01065_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[94][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10637_ (.D(_01066_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[94][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10638_ (.D(_01067_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[94][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10639_ (.D(_01068_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[94][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10640_ (.D(_01069_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[95][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10641_ (.D(_01070_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[95][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10642_ (.D(_01071_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[95][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10643_ (.D(_01072_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[95][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10644_ (.D(_01073_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[95][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10645_ (.D(_01074_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[95][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10646_ (.D(_01075_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[95][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10647_ (.D(_01076_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[95][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10648_ (.D(_01077_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[96][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10649_ (.D(_01078_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[96][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10650_ (.D(_01079_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[96][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10651_ (.D(_01080_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[96][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10652_ (.D(_01081_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[96][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10653_ (.D(_01082_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[96][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10654_ (.D(_01083_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[96][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10655_ (.D(_01084_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[96][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10656_ (.D(_01085_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.bufreg.i_sh_signed ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10657_ (.D(_01086_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.genblk1.align.ctrl_misal ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10658_ (.D(_01087_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[28][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10659_ (.D(_01088_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[28][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10660_ (.D(_01089_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[28][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10661_ (.D(_01090_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[28][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10662_ (.D(_01091_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[28][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10663_ (.D(_01092_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[28][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10664_ (.D(_01093_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[28][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10665_ (.D(_01094_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[28][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10666_ (.D(_01095_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10667_ (.D(_01096_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10668_ (.D(_01097_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10669_ (.D(_01098_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10670_ (.D(_01099_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10671_ (.D(_01100_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10672_ (.D(_01101_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10673_ (.D(_01102_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10674_ (.D(_01103_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10675_ (.D(_01104_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10676_ (.D(_01105_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10677_ (.D(_01106_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10678_ (.D(_01107_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10679_ (.D(_01108_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10680_ (.D(_01109_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10681_ (.D(_01110_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10682_ (.D(_01111_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[101][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10683_ (.D(_01112_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[101][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10684_ (.D(_01113_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[101][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10685_ (.D(_01114_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[101][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10686_ (.D(_01115_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[101][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10687_ (.D(_01116_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[101][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10688_ (.D(_01117_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[101][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10689_ (.D(_01118_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[101][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10690_ (.D(_01119_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[102][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10691_ (.D(_01120_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[102][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10692_ (.D(_01121_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[102][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10693_ (.D(_01122_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[102][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10694_ (.D(_01123_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[102][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10695_ (.D(_01124_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[102][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10696_ (.D(_01125_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[102][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10697_ (.D(_01126_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[102][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10698_ (.D(_01127_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[103][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10699_ (.D(_01128_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[103][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10700_ (.D(_01129_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[103][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10701_ (.D(_01130_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[103][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10702_ (.D(_01131_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[103][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10703_ (.D(_01132_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[103][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10704_ (.D(_01133_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[103][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10705_ (.D(_01134_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[103][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10706_ (.D(_01135_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[104][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10707_ (.D(_01136_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[104][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10708_ (.D(_01137_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[104][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10709_ (.D(_01138_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[104][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10710_ (.D(_01139_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[104][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10711_ (.D(_01140_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[104][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10712_ (.D(_01141_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[104][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10713_ (.D(_01142_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[104][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10714_ (.D(_01143_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[99][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10715_ (.D(_01144_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[99][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10716_ (.D(_01145_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[99][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10717_ (.D(_01146_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[99][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10718_ (.D(_01147_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[99][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10719_ (.D(_01148_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[99][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10720_ (.D(_01149_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[99][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10721_ (.D(_01150_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[99][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10722_ (.D(_01151_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[79][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10723_ (.D(_01152_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[79][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10724_ (.D(_01153_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[79][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10725_ (.D(_01154_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[79][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10726_ (.D(_01155_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[79][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10727_ (.D(_01156_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[79][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10728_ (.D(_01157_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[79][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10729_ (.D(_01158_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[79][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10730_ (.D(_01159_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[105][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10731_ (.D(_01160_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[105][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10732_ (.D(_01161_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[105][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10733_ (.D(_01162_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[105][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10734_ (.D(_01163_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[105][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10735_ (.D(_01164_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[105][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10736_ (.D(_01165_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[105][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10737_ (.D(_01166_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[105][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10738_ (.D(_01167_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[106][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10739_ (.D(_01168_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[106][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10740_ (.D(_01169_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[106][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10741_ (.D(_01170_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[106][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10742_ (.D(_01171_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[106][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10743_ (.D(_01172_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[106][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10744_ (.D(_01173_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[106][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10745_ (.D(_01174_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[106][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10746_ (.D(_01175_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[107][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10747_ (.D(_01176_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[107][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10748_ (.D(_01177_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[107][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10749_ (.D(_01178_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[107][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10750_ (.D(_01179_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[107][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10751_ (.D(_01180_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[107][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10752_ (.D(_01181_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[107][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10753_ (.D(_01182_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[107][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10754_ (.D(_01183_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[83][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10755_ (.D(_01184_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[83][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10756_ (.D(_01185_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[83][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10757_ (.D(_01186_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[83][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10758_ (.D(_01187_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[83][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10759_ (.D(_01188_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[83][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10760_ (.D(_01189_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[83][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10761_ (.D(_01190_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[83][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10762_ (.D(_01191_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[108][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10763_ (.D(_01192_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[108][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10764_ (.D(_01193_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[108][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10765_ (.D(_01194_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[108][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10766_ (.D(_01195_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[108][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10767_ (.D(_01196_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[108][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10768_ (.D(_01197_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[108][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10769_ (.D(_01198_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[108][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10770_ (.D(_01199_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[69][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10771_ (.D(_01200_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[69][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10772_ (.D(_01201_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[69][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10773_ (.D(_01202_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[69][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10774_ (.D(_01203_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[69][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10775_ (.D(_01204_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[69][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10776_ (.D(_01205_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[69][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10777_ (.D(_01206_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[69][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10778_ (.D(_01207_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[84][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10779_ (.D(_01208_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[84][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10780_ (.D(_01209_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[84][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10781_ (.D(_01210_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[84][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10782_ (.D(_01211_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[84][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10783_ (.D(_01212_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[84][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10784_ (.D(_01213_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[84][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10785_ (.D(_01214_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[84][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10786_ (.D(_01215_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[59][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10787_ (.D(_01216_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[59][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10788_ (.D(_01217_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[59][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10789_ (.D(_01218_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[59][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10790_ (.D(_01219_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[59][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10791_ (.D(_01220_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[59][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10792_ (.D(_01221_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[59][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10793_ (.D(_01222_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[59][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10794_ (.D(_01223_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[10][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10795_ (.D(_01224_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[10][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10796_ (.D(_01225_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[10][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10797_ (.D(_01226_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[10][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10798_ (.D(_01227_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[10][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10799_ (.D(_01228_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[10][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10800_ (.D(_01229_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[10][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10801_ (.D(_01230_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[10][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10802_ (.D(_01231_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[85][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10803_ (.D(_01232_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[85][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10804_ (.D(_01233_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[85][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10805_ (.D(_01234_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[85][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10806_ (.D(_01235_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[85][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10807_ (.D(_01236_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[85][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10808_ (.D(_01237_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[85][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10809_ (.D(_01238_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[85][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10810_ (.D(_01239_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[110][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10811_ (.D(_01240_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[110][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10812_ (.D(_01241_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[110][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10813_ (.D(_01242_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[110][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10814_ (.D(_01243_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[110][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10815_ (.D(_01244_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[110][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10816_ (.D(_01245_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[110][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10817_ (.D(_01246_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[110][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10818_ (.D(_01247_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[86][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10819_ (.D(_01248_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[86][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10820_ (.D(_01249_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[86][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10821_ (.D(_01250_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[86][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10822_ (.D(_01251_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[86][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10823_ (.D(_01252_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[86][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10824_ (.D(_01253_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[86][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10825_ (.D(_01254_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[86][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10826_ (.D(_01255_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[111][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10827_ (.D(_01256_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[111][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10828_ (.D(_01257_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[111][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10829_ (.D(_01258_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[111][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10830_ (.D(_01259_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[111][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10831_ (.D(_01260_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[111][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10832_ (.D(_01261_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[111][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10833_ (.D(_01262_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[111][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10834_ (.D(_01263_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[87][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10835_ (.D(_01264_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[87][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10836_ (.D(_01265_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[87][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10837_ (.D(_01266_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[87][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10838_ (.D(_01267_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[87][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10839_ (.D(_01268_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[87][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10840_ (.D(_01269_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[87][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10841_ (.D(_01270_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[87][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10842_ (.D(_01271_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[88][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10843_ (.D(_01272_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[88][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10844_ (.D(_01273_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[88][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10845_ (.D(_01274_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[88][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10846_ (.D(_01275_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[88][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10847_ (.D(_01276_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[88][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10848_ (.D(_01277_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[88][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10849_ (.D(_01278_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[88][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10850_ (.D(_01279_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.genblk3.csr.mcause3_0[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10851_ (.D(_01280_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.genblk3.csr.mcause3_0[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10852_ (.D(_01281_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.genblk3.csr.mcause3_0[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10853_ (.D(_01282_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.genblk3.csr.mcause3_0[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10854_ (.D(_01283_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.genblk3.csr.mcause31 ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10855_ (.D(_01284_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.genblk3.csr.mstatus_mpie ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10856_ (.D(_01285_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.genblk3.csr.mie_mtie ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10857_ (.D(_01286_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.genblk3.csr.mstatus_mie ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10858_ (.D(_01287_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.ctrl.i_iscomp ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10859_ (.D(_01288_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.genblk3.csr.o_new_irq ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10860_ (.D(_01289_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[27][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10861_ (.D(_01290_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[27][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10862_ (.D(_01291_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[27][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10863_ (.D(_01292_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[27][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10864_ (.D(_01293_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[27][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10865_ (.D(_01294_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[27][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10866_ (.D(_01295_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[27][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10867_ (.D(_01296_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[27][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10868_ (.D(_01297_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[26][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10869_ (.D(_01298_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[26][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10870_ (.D(_01299_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[26][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10871_ (.D(_01300_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[26][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10872_ (.D(_01301_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[26][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10873_ (.D(_01302_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[26][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10874_ (.D(_01303_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[26][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10875_ (.D(_01304_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[26][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10876_ (.D(_01305_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[25][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10877_ (.D(_01306_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[25][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10878_ (.D(_01307_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[25][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10879_ (.D(_01308_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[25][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10880_ (.D(_01309_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[25][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10881_ (.D(_01310_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[25][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10882_ (.D(_01311_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[25][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10883_ (.D(_01312_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[25][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10884_ (.D(_01313_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[24][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10885_ (.D(_01314_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[24][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10886_ (.D(_01315_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[24][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10887_ (.D(_01316_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[24][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10888_ (.D(_01317_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[24][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10889_ (.D(_01318_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[24][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10890_ (.D(_01319_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[24][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10891_ (.D(_01320_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[24][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10892_ (.D(_01321_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[0][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10893_ (.D(_01322_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[0][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10894_ (.D(_01323_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[0][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10895_ (.D(_01324_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[0][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10896_ (.D(_01325_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[0][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10897_ (.D(_01326_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[0][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10898_ (.D(_01327_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[0][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10899_ (.D(_01328_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[0][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10900_ (.D(_01329_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[98][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10901_ (.D(_01330_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[98][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10902_ (.D(_01331_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[98][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10903_ (.D(_01332_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[98][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10904_ (.D(_01333_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[98][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10905_ (.D(_01334_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[98][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10906_ (.D(_01335_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[98][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10907_ (.D(_01336_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[98][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10908_ (.D(_01337_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[100][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10909_ (.D(_01338_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[100][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10910_ (.D(_01339_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[100][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10911_ (.D(_01340_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[100][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10912_ (.D(_01341_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[100][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10913_ (.D(_01342_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[100][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10914_ (.D(_01343_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[100][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10915_ (.D(_01344_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[100][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10916_ (.D(_01345_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[89][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10917_ (.D(_01346_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[89][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10918_ (.D(_01347_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[89][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10919_ (.D(_01348_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[89][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10920_ (.D(_01349_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[89][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10921_ (.D(_01350_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[89][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10922_ (.D(_01351_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[89][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10923_ (.D(_01352_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[89][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10924_ (.D(_00025_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.regzero ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10925_ (.D(_01353_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[23][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10926_ (.D(_01354_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[23][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10927_ (.D(_01355_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[23][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10928_ (.D(_01356_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[23][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10929_ (.D(_01357_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[23][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10930_ (.D(_01358_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[23][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10931_ (.D(_01359_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[23][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10932_ (.D(_01360_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram.memory[23][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10933_ (.D(_01361_),
    .CLK(io_in[4]),
    .Q(\u_cpu.cpu.state.ibus_cyc ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10934_ (.D(\u_cpu.rf_ram_if.wdata0_r[1] ),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram_if.wdata0_r[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10935_ (.D(\u_cpu.rf_ram_if.wdata0_r[2] ),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram_if.wdata0_r[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10936_ (.D(\u_cpu.rf_ram_if.wdata0_r[3] ),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram_if.wdata0_r[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10937_ (.D(\u_cpu.rf_ram_if.wdata0_r[4] ),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram_if.wdata0_r[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10938_ (.D(\u_cpu.rf_ram_if.wdata0_r[5] ),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram_if.wdata0_r[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10939_ (.D(\u_cpu.rf_ram_if.wdata0_r[6] ),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram_if.wdata0_r[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10940_ (.D(\u_cpu.cpu.o_wdata0 ),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram_if.wdata0_r[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10941_ (.D(\u_cpu.rf_ram_if.wtrig0 ),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram_if.genblk1.wtrig0_r ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10942_ (.D(_01362_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram_if.rdata1[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10943_ (.D(_01363_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram_if.rdata0[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10944_ (.D(_01364_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram_if.rgnt ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10945_ (.D(\u_cpu.rf_ram_if.rtrig0 ),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram_if.rtrig1 ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10946_ (.D(_01365_),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram_if.rcnt[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10947_ (.D(\u_cpu.rf_ram_if.wdata1_r[1] ),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram_if.wdata1_r[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10948_ (.D(\u_cpu.rf_ram_if.wdata1_r[2] ),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram_if.wdata1_r[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10949_ (.D(\u_cpu.rf_ram_if.wdata1_r[3] ),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram_if.wdata1_r[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10950_ (.D(\u_cpu.rf_ram_if.wdata1_r[4] ),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram_if.wdata1_r[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10951_ (.D(\u_cpu.rf_ram_if.wdata1_r[5] ),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram_if.wdata1_r[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10952_ (.D(\u_cpu.rf_ram_if.wdata1_r[6] ),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram_if.wdata1_r[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10953_ (.D(\u_cpu.rf_ram_if.wdata1_r[7] ),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram_if.wdata1_r[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10954_ (.D(\u_cpu.cpu.o_wdata1 ),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram_if.wdata1_r[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10955_ (.D(\u_cpu.cpu.o_wen0 ),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram_if.wen0_r ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10956_ (.D(\u_cpu.cpu.o_wen1 ),
    .CLK(io_in[4]),
    .Q(\u_cpu.rf_ram_if.wen1_r ));
 gf180mcu_fd_sc_mcu7t5v0__tieh _10957_ (.Z(_04690_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _10958_ (.Z(_04691_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _10959_ (.Z(_04692_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _10960_ (.Z(_04693_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _10961_ (.Z(_04694_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _10962_ (.Z(_04695_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _10963_ (.Z(_04696_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _10964_ (.Z(_04697_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _10965_ (.Z(_04698_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _10966_ (.Z(_04699_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _10967_ (.Z(_04700_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _10968_ (.Z(_04701_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _10969_ (.Z(_04702_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _10970_ (.Z(_04703_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _10971_ (.Z(_04704_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _10972_ (.Z(_04705_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _10973_ (.Z(_04706_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _10974_ (.Z(_04707_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _10975_ (.Z(_04708_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _10976_ (.Z(_04709_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _10977_ (.Z(_04710_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _10978_ (.Z(_04711_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _10979_ (.Z(_04712_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _10980_ (.Z(_04713_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _10981_ (.Z(_04714_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _10982_ (.Z(_04715_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _10983_ (.Z(_04716_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _10984_ (.Z(_04717_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _10985_ (.Z(_04718_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _10986_ (.Z(_04719_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _10987_ (.Z(_04720_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _10988_ (.Z(_04721_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _10989_ (.Z(_04722_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _10990_ (.Z(_04723_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _10991_ (.Z(_04724_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _10992_ (.Z(_04725_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _10993_ (.Z(_04726_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _10994_ (.Z(_04727_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _10995_ (.Z(_04728_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _10996_ (.Z(_04729_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _10997_ (.Z(_04730_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _10998_ (.Z(_04731_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _10999_ (.Z(_04732_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _11000_ (.Z(_04733_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _11001_ (.Z(_04734_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _11002_ (.Z(_04735_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _11003_ (.Z(_04736_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _11004_ (.Z(_04737_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _11005_ (.Z(_04738_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _11006_ (.Z(_04739_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _11007_ (.Z(_04740_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _11008_ (.Z(_04741_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _11009_ (.Z(_04742_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _11010_ (.Z(_04743_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _11011_ (.Z(_04744_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _11012_ (.Z(_04745_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _11013_ (.Z(_04746_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _11014_ (.Z(_04747_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _11015_ (.Z(_04748_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _11016_ (.Z(_04749_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _11017_ (.Z(_04750_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _11018_ (.Z(_04751_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _11019_ (.Z(_04752_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _11020_ (.Z(_04753_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _11021_ (.Z(_04754_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _11022_ (.Z(_04755_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _11023_ (.Z(_04756_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _11024_ (.Z(_04757_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _11025_ (.Z(_04758_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _11026_ (.Z(_04759_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _11027_ (.Z(_04760_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _11028_ (.Z(_04761_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _11029_ (.Z(_04762_));
 gf180mcu_fd_sc_mcu7t5v0__tieh _11030_ (.Z(_04763_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _11031_ (.ZN(_04764_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _11032_ (.ZN(_04765_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _11033_ (.ZN(_04766_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _11034_ (.ZN(_04767_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _11035_ (.ZN(_04768_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _11036_ (.ZN(_04769_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _11037_ (.ZN(_04770_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _11038_ (.ZN(_04771_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _11039_ (.ZN(_04772_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _11040_ (.ZN(_04773_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _11041_ (.ZN(_04774_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _11042_ (.ZN(_04775_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _11043_ (.ZN(_04776_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _11044_ (.ZN(_04777_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _11045_ (.ZN(_04778_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _11046_ (.ZN(_04779_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _11047_ (.ZN(_04780_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _11048_ (.ZN(_04781_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _11049_ (.ZN(_04782_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _11050_ (.ZN(_04783_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _11051_ (.ZN(_04784_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _11052_ (.ZN(_04785_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _11053_ (.ZN(_04786_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _11054_ (.ZN(_04787_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _11055_ (.ZN(_04788_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _11056_ (.ZN(_04789_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _11057_ (.ZN(_04790_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _11058_ (.ZN(_04791_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _11059_ (.ZN(_04792_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _11060_ (.ZN(_04793_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _11061_ (.ZN(_04794_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _11062_ (.ZN(_04795_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _11063_ (.ZN(_04796_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _11064_ (.ZN(_04797_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _11065_ (.ZN(_04798_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _11066_ (.ZN(_04799_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _11067_ (.ZN(_04800_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _11068_ (.ZN(_04801_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _11069_ (.ZN(_04802_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _11070_ (.ZN(_04803_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _11071_ (.ZN(_04804_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _11072_ (.ZN(_04805_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _11073_ (.ZN(_04806_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _11074_ (.ZN(_04807_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _11075_ (.ZN(_04808_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _11076_ (.ZN(_04809_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _11077_ (.ZN(_04810_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _11078_ (.ZN(_04811_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _11079_ (.ZN(_04812_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _11080_ (.ZN(_04813_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _11081_ (.ZN(_04814_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _11082_ (.ZN(_04815_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _11083_ (.ZN(_04816_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _11084_ (.ZN(_04817_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _11085_ (.ZN(_04818_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _11086_ (.ZN(_04819_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _11087_ (.ZN(_04820_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _11088_ (.ZN(_04821_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _11089_ (.ZN(_04822_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _11090_ (.ZN(_04823_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _11091_ (.ZN(_04824_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _11092_ (.ZN(_04825_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _11093_ (.ZN(_04826_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _11094_ (.ZN(_04827_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _11095_ (.ZN(_04828_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _11096_ (.ZN(_04829_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _11097_ (.ZN(_04830_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _11098_ (.ZN(_04831_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _11099_ (.ZN(_04832_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _11100_ (.ZN(_04833_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _11101_ (.ZN(_04834_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _11102_ (.ZN(_04835_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _11103_ (.ZN(_04836_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _11104_ (.ZN(_04837_));
 gf180mcu_fd_sc_mcu7t5v0__tiel _11105_ (.ZN(io_oeb[0]));
 gf180mcu_fd_sc_mcu7t5v0__tiel _11106_ (.ZN(io_oeb[1]));
 gf180mcu_fd_sc_mcu7t5v0__tiel _11107_ (.ZN(io_oeb[2]));
 gf180mcu_fd_sc_mcu7t5v0__tiel _11108_ (.ZN(io_oeb[3]));
 gf180mcu_fd_sc_mcu7t5v0__tiel _11109_ (.ZN(io_oeb[4]));
 gf180mcu_fd_sc_mcu7t5v0__tiel _11110_ (.ZN(io_out[2]));
 gf180mcu_fd_sc_mcu7t5v0__tiel _11111_ (.ZN(io_out[3]));
 gf180mcu_fd_sc_mcu7t5v0__tiel _11112_ (.ZN(io_out[4]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11113_ (.I(\u_scanchain_local.clk_out ),
    .Z(io_out[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11114_ (.I(\u_scanchain_local.data_out ),
    .Z(io_out[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 \u_scanchain_local.input_buf_clk  (.I(io_in[0]),
    .Z(\u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__dffnq_1 \u_scanchain_local.out_flop  (.D(\u_scanchain_local.module_data_in[69] ),
    .CLKN(\u_scanchain_local.clk ),
    .Q(\u_scanchain_local.data_out_i ));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 \u_scanchain_local.output_buffers[2]  (.I(\u_scanchain_local.data_out_i ),
    .Z(\u_scanchain_local.data_out ));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 \u_scanchain_local.output_buffers[3]  (.I(\u_scanchain_local.clk ),
    .Z(\u_scanchain_local.clk_out ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[0]  (.D(io_in[2]),
    .SE(io_in[3]),
    .SI(\u_arbiter.o_wb_cpu_cyc ),
    .CLK(\u_scanchain_local.clk ),
    .Q(\u_cpu.cpu.genblk3.csr.i_mtip ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[10]  (.D(\u_arbiter.i_wb_cpu_rdt[7] ),
    .SE(io_in[3]),
    .SI(\u_arbiter.i_wb_cpu_dbus_dat[4] ),
    .CLK(\u_scanchain_local.clk ),
    .Q(\u_arbiter.i_wb_cpu_rdt[8] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[11]  (.D(\u_arbiter.i_wb_cpu_rdt[8] ),
    .SE(io_in[3]),
    .SI(\u_arbiter.i_wb_cpu_dbus_dat[5] ),
    .CLK(\u_scanchain_local.clk ),
    .Q(\u_arbiter.i_wb_cpu_rdt[9] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[12]  (.D(\u_arbiter.i_wb_cpu_rdt[9] ),
    .SE(io_in[3]),
    .SI(\u_arbiter.i_wb_cpu_dbus_dat[6] ),
    .CLK(\u_scanchain_local.clk ),
    .Q(\u_arbiter.i_wb_cpu_rdt[10] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[13]  (.D(\u_arbiter.i_wb_cpu_rdt[10] ),
    .SE(io_in[3]),
    .SI(\u_arbiter.i_wb_cpu_dbus_dat[7] ),
    .CLK(\u_scanchain_local.clk ),
    .Q(\u_arbiter.i_wb_cpu_rdt[11] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[14]  (.D(\u_arbiter.i_wb_cpu_rdt[11] ),
    .SE(io_in[3]),
    .SI(\u_arbiter.i_wb_cpu_dbus_dat[8] ),
    .CLK(\u_scanchain_local.clk ),
    .Q(\u_arbiter.i_wb_cpu_rdt[12] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[15]  (.D(\u_arbiter.i_wb_cpu_rdt[12] ),
    .SE(io_in[3]),
    .SI(\u_arbiter.i_wb_cpu_dbus_dat[9] ),
    .CLK(\u_scanchain_local.clk ),
    .Q(\u_arbiter.i_wb_cpu_rdt[13] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[16]  (.D(\u_arbiter.i_wb_cpu_rdt[13] ),
    .SE(io_in[3]),
    .SI(\u_arbiter.i_wb_cpu_dbus_dat[10] ),
    .CLK(\u_scanchain_local.clk ),
    .Q(\u_arbiter.i_wb_cpu_rdt[14] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[17]  (.D(\u_arbiter.i_wb_cpu_rdt[14] ),
    .SE(io_in[3]),
    .SI(\u_arbiter.i_wb_cpu_dbus_dat[11] ),
    .CLK(\u_scanchain_local.clk ),
    .Q(\u_arbiter.i_wb_cpu_rdt[15] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[18]  (.D(\u_arbiter.i_wb_cpu_rdt[15] ),
    .SE(io_in[3]),
    .SI(\u_arbiter.i_wb_cpu_dbus_dat[12] ),
    .CLK(\u_scanchain_local.clk ),
    .Q(\u_arbiter.i_wb_cpu_rdt[16] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[19]  (.D(\u_arbiter.i_wb_cpu_rdt[16] ),
    .SE(io_in[3]),
    .SI(\u_arbiter.i_wb_cpu_dbus_dat[13] ),
    .CLK(\u_scanchain_local.clk ),
    .Q(\u_arbiter.i_wb_cpu_rdt[17] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[1]  (.D(\u_cpu.cpu.genblk3.csr.i_mtip ),
    .SE(io_in[3]),
    .SI(\u_arbiter.o_wb_cpu_we ),
    .CLK(\u_scanchain_local.clk ),
    .Q(\u_arbiter.i_wb_cpu_ack ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[20]  (.D(\u_arbiter.i_wb_cpu_rdt[17] ),
    .SE(io_in[3]),
    .SI(\u_arbiter.i_wb_cpu_dbus_dat[14] ),
    .CLK(\u_scanchain_local.clk ),
    .Q(\u_arbiter.i_wb_cpu_rdt[18] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[21]  (.D(\u_arbiter.i_wb_cpu_rdt[18] ),
    .SE(io_in[3]),
    .SI(\u_arbiter.i_wb_cpu_dbus_dat[15] ),
    .CLK(\u_scanchain_local.clk ),
    .Q(\u_arbiter.i_wb_cpu_rdt[19] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[22]  (.D(\u_arbiter.i_wb_cpu_rdt[19] ),
    .SE(io_in[3]),
    .SI(\u_arbiter.i_wb_cpu_dbus_dat[16] ),
    .CLK(\u_scanchain_local.clk ),
    .Q(\u_arbiter.i_wb_cpu_rdt[20] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[23]  (.D(\u_arbiter.i_wb_cpu_rdt[20] ),
    .SE(io_in[3]),
    .SI(\u_arbiter.i_wb_cpu_dbus_dat[17] ),
    .CLK(\u_scanchain_local.clk ),
    .Q(\u_arbiter.i_wb_cpu_rdt[21] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[24]  (.D(\u_arbiter.i_wb_cpu_rdt[21] ),
    .SE(io_in[3]),
    .SI(\u_arbiter.i_wb_cpu_dbus_dat[18] ),
    .CLK(\u_scanchain_local.clk ),
    .Q(\u_arbiter.i_wb_cpu_rdt[22] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[25]  (.D(\u_arbiter.i_wb_cpu_rdt[22] ),
    .SE(io_in[3]),
    .SI(\u_arbiter.i_wb_cpu_dbus_dat[19] ),
    .CLK(\u_scanchain_local.clk ),
    .Q(\u_arbiter.i_wb_cpu_rdt[23] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[26]  (.D(\u_arbiter.i_wb_cpu_rdt[23] ),
    .SE(io_in[3]),
    .SI(\u_arbiter.i_wb_cpu_dbus_dat[20] ),
    .CLK(\u_scanchain_local.clk ),
    .Q(\u_arbiter.i_wb_cpu_rdt[24] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[27]  (.D(\u_arbiter.i_wb_cpu_rdt[24] ),
    .SE(io_in[3]),
    .SI(\u_arbiter.i_wb_cpu_dbus_dat[21] ),
    .CLK(\u_scanchain_local.clk ),
    .Q(\u_arbiter.i_wb_cpu_rdt[25] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[28]  (.D(\u_arbiter.i_wb_cpu_rdt[25] ),
    .SE(io_in[3]),
    .SI(\u_arbiter.i_wb_cpu_dbus_dat[22] ),
    .CLK(\u_scanchain_local.clk ),
    .Q(\u_arbiter.i_wb_cpu_rdt[26] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[29]  (.D(\u_arbiter.i_wb_cpu_rdt[26] ),
    .SE(io_in[3]),
    .SI(\u_arbiter.i_wb_cpu_dbus_dat[23] ),
    .CLK(\u_scanchain_local.clk ),
    .Q(\u_arbiter.i_wb_cpu_rdt[27] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[2]  (.D(\u_arbiter.i_wb_cpu_ack ),
    .SE(io_in[3]),
    .SI(\u_arbiter.i_wb_cpu_dbus_sel[0] ),
    .CLK(\u_scanchain_local.clk ),
    .Q(\u_arbiter.i_wb_cpu_rdt[0] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[30]  (.D(\u_arbiter.i_wb_cpu_rdt[27] ),
    .SE(io_in[3]),
    .SI(\u_arbiter.i_wb_cpu_dbus_dat[24] ),
    .CLK(\u_scanchain_local.clk ),
    .Q(\u_arbiter.i_wb_cpu_rdt[28] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[31]  (.D(\u_arbiter.i_wb_cpu_rdt[28] ),
    .SE(io_in[3]),
    .SI(\u_arbiter.i_wb_cpu_dbus_dat[25] ),
    .CLK(\u_scanchain_local.clk ),
    .Q(\u_arbiter.i_wb_cpu_rdt[29] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[32]  (.D(\u_arbiter.i_wb_cpu_rdt[29] ),
    .SE(io_in[3]),
    .SI(\u_arbiter.i_wb_cpu_dbus_dat[26] ),
    .CLK(\u_scanchain_local.clk ),
    .Q(\u_arbiter.i_wb_cpu_rdt[30] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[33]  (.D(\u_arbiter.i_wb_cpu_rdt[30] ),
    .SE(io_in[3]),
    .SI(\u_arbiter.i_wb_cpu_dbus_dat[27] ),
    .CLK(\u_scanchain_local.clk ),
    .Q(\u_arbiter.i_wb_cpu_rdt[31] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[34]  (.D(\u_arbiter.i_wb_cpu_rdt[31] ),
    .SE(io_in[3]),
    .SI(\u_arbiter.i_wb_cpu_dbus_dat[28] ),
    .CLK(\u_scanchain_local.clk ),
    .Q(\u_scanchain_local.module_data_in[34] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[35]  (.D(\u_scanchain_local.module_data_in[34] ),
    .SE(io_in[3]),
    .SI(\u_arbiter.i_wb_cpu_dbus_dat[29] ),
    .CLK(\u_scanchain_local.clk ),
    .Q(\u_scanchain_local.module_data_in[35] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[36]  (.D(\u_scanchain_local.module_data_in[35] ),
    .SE(io_in[3]),
    .SI(\u_arbiter.i_wb_cpu_dbus_dat[30] ),
    .CLK(\u_scanchain_local.clk ),
    .Q(\u_scanchain_local.module_data_in[36] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[37]  (.D(\u_scanchain_local.module_data_in[36] ),
    .SE(io_in[3]),
    .SI(\u_arbiter.i_wb_cpu_dbus_dat[31] ),
    .CLK(\u_scanchain_local.clk ),
    .Q(\u_scanchain_local.module_data_in[37] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[38]  (.D(\u_scanchain_local.module_data_in[37] ),
    .SE(io_in[3]),
    .SI(\u_arbiter.o_wb_cpu_adr[0] ),
    .CLK(\u_scanchain_local.clk ),
    .Q(\u_scanchain_local.module_data_in[38] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[39]  (.D(\u_scanchain_local.module_data_in[38] ),
    .SE(io_in[3]),
    .SI(\u_arbiter.o_wb_cpu_adr[1] ),
    .CLK(\u_scanchain_local.clk ),
    .Q(\u_scanchain_local.module_data_in[39] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[3]  (.D(\u_arbiter.i_wb_cpu_rdt[0] ),
    .SE(io_in[3]),
    .SI(\u_arbiter.i_wb_cpu_dbus_sel[1] ),
    .CLK(\u_scanchain_local.clk ),
    .Q(\u_arbiter.i_wb_cpu_rdt[1] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[40]  (.D(\u_scanchain_local.module_data_in[39] ),
    .SE(io_in[3]),
    .SI(\u_arbiter.o_wb_cpu_adr[2] ),
    .CLK(\u_scanchain_local.clk ),
    .Q(\u_scanchain_local.module_data_in[40] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[41]  (.D(\u_scanchain_local.module_data_in[40] ),
    .SE(io_in[3]),
    .SI(\u_arbiter.o_wb_cpu_adr[3] ),
    .CLK(\u_scanchain_local.clk ),
    .Q(\u_scanchain_local.module_data_in[41] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[42]  (.D(\u_scanchain_local.module_data_in[41] ),
    .SE(io_in[3]),
    .SI(\u_arbiter.o_wb_cpu_adr[4] ),
    .CLK(\u_scanchain_local.clk ),
    .Q(\u_scanchain_local.module_data_in[42] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[43]  (.D(\u_scanchain_local.module_data_in[42] ),
    .SE(io_in[3]),
    .SI(\u_arbiter.o_wb_cpu_adr[5] ),
    .CLK(\u_scanchain_local.clk ),
    .Q(\u_scanchain_local.module_data_in[43] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[44]  (.D(\u_scanchain_local.module_data_in[43] ),
    .SE(io_in[3]),
    .SI(\u_arbiter.o_wb_cpu_adr[6] ),
    .CLK(\u_scanchain_local.clk ),
    .Q(\u_scanchain_local.module_data_in[44] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[45]  (.D(\u_scanchain_local.module_data_in[44] ),
    .SE(io_in[3]),
    .SI(\u_arbiter.o_wb_cpu_adr[7] ),
    .CLK(\u_scanchain_local.clk ),
    .Q(\u_scanchain_local.module_data_in[45] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[46]  (.D(\u_scanchain_local.module_data_in[45] ),
    .SE(io_in[3]),
    .SI(\u_arbiter.o_wb_cpu_adr[8] ),
    .CLK(\u_scanchain_local.clk ),
    .Q(\u_scanchain_local.module_data_in[46] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[47]  (.D(\u_scanchain_local.module_data_in[46] ),
    .SE(io_in[3]),
    .SI(\u_arbiter.o_wb_cpu_adr[9] ),
    .CLK(\u_scanchain_local.clk ),
    .Q(\u_scanchain_local.module_data_in[47] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[48]  (.D(\u_scanchain_local.module_data_in[47] ),
    .SE(io_in[3]),
    .SI(\u_arbiter.o_wb_cpu_adr[10] ),
    .CLK(\u_scanchain_local.clk ),
    .Q(\u_scanchain_local.module_data_in[48] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[49]  (.D(\u_scanchain_local.module_data_in[48] ),
    .SE(io_in[3]),
    .SI(\u_arbiter.o_wb_cpu_adr[11] ),
    .CLK(\u_scanchain_local.clk ),
    .Q(\u_scanchain_local.module_data_in[49] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[4]  (.D(\u_arbiter.i_wb_cpu_rdt[1] ),
    .SE(io_in[3]),
    .SI(\u_arbiter.i_wb_cpu_dbus_sel[2] ),
    .CLK(\u_scanchain_local.clk ),
    .Q(\u_arbiter.i_wb_cpu_rdt[2] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[50]  (.D(\u_scanchain_local.module_data_in[49] ),
    .SE(io_in[3]),
    .SI(\u_arbiter.o_wb_cpu_adr[12] ),
    .CLK(\u_scanchain_local.clk ),
    .Q(\u_scanchain_local.module_data_in[50] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[51]  (.D(\u_scanchain_local.module_data_in[50] ),
    .SE(io_in[3]),
    .SI(\u_arbiter.o_wb_cpu_adr[13] ),
    .CLK(\u_scanchain_local.clk ),
    .Q(\u_scanchain_local.module_data_in[51] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[52]  (.D(\u_scanchain_local.module_data_in[51] ),
    .SE(io_in[3]),
    .SI(\u_arbiter.o_wb_cpu_adr[14] ),
    .CLK(\u_scanchain_local.clk ),
    .Q(\u_scanchain_local.module_data_in[52] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[53]  (.D(\u_scanchain_local.module_data_in[52] ),
    .SE(io_in[3]),
    .SI(\u_arbiter.o_wb_cpu_adr[15] ),
    .CLK(\u_scanchain_local.clk ),
    .Q(\u_scanchain_local.module_data_in[53] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[54]  (.D(\u_scanchain_local.module_data_in[53] ),
    .SE(io_in[3]),
    .SI(\u_arbiter.o_wb_cpu_adr[16] ),
    .CLK(\u_scanchain_local.clk ),
    .Q(\u_scanchain_local.module_data_in[54] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[55]  (.D(\u_scanchain_local.module_data_in[54] ),
    .SE(io_in[3]),
    .SI(\u_arbiter.o_wb_cpu_adr[17] ),
    .CLK(\u_scanchain_local.clk ),
    .Q(\u_scanchain_local.module_data_in[55] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[56]  (.D(\u_scanchain_local.module_data_in[55] ),
    .SE(io_in[3]),
    .SI(\u_arbiter.o_wb_cpu_adr[18] ),
    .CLK(\u_scanchain_local.clk ),
    .Q(\u_scanchain_local.module_data_in[56] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[57]  (.D(\u_scanchain_local.module_data_in[56] ),
    .SE(io_in[3]),
    .SI(\u_arbiter.o_wb_cpu_adr[19] ),
    .CLK(\u_scanchain_local.clk ),
    .Q(\u_scanchain_local.module_data_in[57] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[58]  (.D(\u_scanchain_local.module_data_in[57] ),
    .SE(io_in[3]),
    .SI(\u_arbiter.o_wb_cpu_adr[20] ),
    .CLK(\u_scanchain_local.clk ),
    .Q(\u_scanchain_local.module_data_in[58] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[59]  (.D(\u_scanchain_local.module_data_in[58] ),
    .SE(io_in[3]),
    .SI(\u_arbiter.o_wb_cpu_adr[21] ),
    .CLK(\u_scanchain_local.clk ),
    .Q(\u_scanchain_local.module_data_in[59] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[5]  (.D(\u_arbiter.i_wb_cpu_rdt[2] ),
    .SE(io_in[3]),
    .SI(\u_arbiter.i_wb_cpu_dbus_sel[3] ),
    .CLK(\u_scanchain_local.clk ),
    .Q(\u_arbiter.i_wb_cpu_rdt[3] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[60]  (.D(\u_scanchain_local.module_data_in[59] ),
    .SE(io_in[3]),
    .SI(\u_arbiter.o_wb_cpu_adr[22] ),
    .CLK(\u_scanchain_local.clk ),
    .Q(\u_scanchain_local.module_data_in[60] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[61]  (.D(\u_scanchain_local.module_data_in[60] ),
    .SE(io_in[3]),
    .SI(\u_arbiter.o_wb_cpu_adr[23] ),
    .CLK(\u_scanchain_local.clk ),
    .Q(\u_scanchain_local.module_data_in[61] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[62]  (.D(\u_scanchain_local.module_data_in[61] ),
    .SE(io_in[3]),
    .SI(\u_arbiter.o_wb_cpu_adr[24] ),
    .CLK(\u_scanchain_local.clk ),
    .Q(\u_scanchain_local.module_data_in[62] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[63]  (.D(\u_scanchain_local.module_data_in[62] ),
    .SE(io_in[3]),
    .SI(\u_arbiter.o_wb_cpu_adr[25] ),
    .CLK(\u_scanchain_local.clk ),
    .Q(\u_scanchain_local.module_data_in[63] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[64]  (.D(\u_scanchain_local.module_data_in[63] ),
    .SE(io_in[3]),
    .SI(\u_arbiter.o_wb_cpu_adr[26] ),
    .CLK(\u_scanchain_local.clk ),
    .Q(\u_scanchain_local.module_data_in[64] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[65]  (.D(\u_scanchain_local.module_data_in[64] ),
    .SE(io_in[3]),
    .SI(\u_arbiter.o_wb_cpu_adr[27] ),
    .CLK(\u_scanchain_local.clk ),
    .Q(\u_scanchain_local.module_data_in[65] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[66]  (.D(\u_scanchain_local.module_data_in[65] ),
    .SE(io_in[3]),
    .SI(\u_arbiter.o_wb_cpu_adr[28] ),
    .CLK(\u_scanchain_local.clk ),
    .Q(\u_scanchain_local.module_data_in[66] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[67]  (.D(\u_scanchain_local.module_data_in[66] ),
    .SE(io_in[3]),
    .SI(\u_arbiter.o_wb_cpu_adr[29] ),
    .CLK(\u_scanchain_local.clk ),
    .Q(\u_scanchain_local.module_data_in[67] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[68]  (.D(\u_scanchain_local.module_data_in[67] ),
    .SE(io_in[3]),
    .SI(\u_arbiter.o_wb_cpu_adr[30] ),
    .CLK(\u_scanchain_local.clk ),
    .Q(\u_scanchain_local.module_data_in[68] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[69]  (.D(\u_scanchain_local.module_data_in[68] ),
    .SE(io_in[3]),
    .SI(\u_arbiter.o_wb_cpu_adr[31] ),
    .CLK(\u_scanchain_local.clk ),
    .Q(\u_scanchain_local.module_data_in[69] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[6]  (.D(\u_arbiter.i_wb_cpu_rdt[3] ),
    .SE(io_in[3]),
    .SI(\u_arbiter.i_wb_cpu_dbus_dat[0] ),
    .CLK(\u_scanchain_local.clk ),
    .Q(\u_arbiter.i_wb_cpu_rdt[4] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[7]  (.D(\u_arbiter.i_wb_cpu_rdt[4] ),
    .SE(io_in[3]),
    .SI(\u_arbiter.i_wb_cpu_dbus_dat[1] ),
    .CLK(\u_scanchain_local.clk ),
    .Q(\u_arbiter.i_wb_cpu_rdt[5] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[8]  (.D(\u_arbiter.i_wb_cpu_rdt[5] ),
    .SE(io_in[3]),
    .SI(\u_arbiter.i_wb_cpu_dbus_dat[2] ),
    .CLK(\u_scanchain_local.clk ),
    .Q(\u_arbiter.i_wb_cpu_rdt[6] ));
 gf180mcu_fd_sc_mcu7t5v0__sdffq_1 \u_scanchain_local.scan_flop[9]  (.D(\u_arbiter.i_wb_cpu_rdt[6] ),
    .SE(io_in[3]),
    .SI(\u_arbiter.i_wb_cpu_dbus_dat[3] ),
    .CLK(\u_scanchain_local.clk ),
    .Q(\u_arbiter.i_wb_cpu_rdt[7] ));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_0 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_6 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_7 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_8 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_9 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_10 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_11 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_12 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_13 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_14 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_15 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_16 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_17 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_18 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_19 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_20 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_21 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_22 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_23 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_24 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_25 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_26 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_27 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_28 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_29 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_30 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_31 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_32 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_33 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_34 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_35 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_36 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_37 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_38 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_39 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_40 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_41 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_42 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_43 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_44 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_45 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_46 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_47 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_48 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_49 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_50 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_51 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_52 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_53 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_54 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_55 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_56 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_57 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_58 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_59 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_60 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_61 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_62 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_63 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_64 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_65 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_66 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_67 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_68 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_69 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_70 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_71 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_72 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_73 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_74 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_75 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_76 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_77 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_78 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_79 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_80 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_81 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_82 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_83 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_84 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_85 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_86 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_87 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_88 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_89 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_90 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_91 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_92 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_93 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_94 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_95 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_96 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_97 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_98 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_99 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_100 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_101 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_102 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_103 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_104 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_105 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_106 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_107 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_108 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_109 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_110 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_111 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_112 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_113 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_114 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_115 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_116 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_117 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_118 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_119 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_120 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_121 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_122 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_123 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_124 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_125 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_126 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_127 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_128 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_129 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_130 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_131 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_132 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_133 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_134 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_135 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_136 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_137 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_138 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_139 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_140 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_141 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_142 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_143 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_144 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_145 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_146 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_147 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_148 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_149 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_150 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_151 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_152 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_153 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_154 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_155 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_156 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_157 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_158 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_159 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_160 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_161 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_162 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_163 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_164 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_165 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_166 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_167 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_168 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_169 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_170 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_171 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_172 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_173 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_174 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_175 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_176 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_177 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_178 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_179 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_180 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_181 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_182 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_183 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_184 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_185 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_186 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_187 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_188 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_189 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_190 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_191 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_192 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_193 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_194 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_195 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_196 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_197 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_198 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_199 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_200 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_201 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_202 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_203 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_204 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_205 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_206 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_207 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_208 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_209 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_210 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_211 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_212 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_213 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_214 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_215 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_216 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_217 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_218 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_219 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_220 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_221 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_222 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_223 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_224 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_225 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_226 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_227 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_228 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_229 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_230 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_231 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_232 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_233 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_234 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_235 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_236 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_237 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_238 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_239 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_240 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_241 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_242 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_243 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_244 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_245 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_246 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_247 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_248 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_249 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_250 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_251 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_252 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_253 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_254 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_255 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_256 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_257 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_258 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_259 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_260 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_261 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_262 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_263 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_264 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_265 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_266 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_267 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_268 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_269 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_270 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_271 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_272 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_273 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_274 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_275 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_276 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_277 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_278 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_279 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_280 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_281 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_282 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_283 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_284 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_285 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_286 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_287 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_288 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2788 ();
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09993__D (.I(_00000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09996__D (.I(_00003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10455__D (.I(_00888_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04897__A2 (.I(_01368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04893__A2 (.I(_01368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04877__I (.I(_01368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04874__A2 (.I(_01368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04869__C (.I(_01368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04841__I (.I(_01368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07738__B (.I(_01369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05907__A1 (.I(_01369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05886__A2 (.I(_01369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05882__A1 (.I(_01369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05875__A1 (.I(_01369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05870__B (.I(_01369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05848__A1 (.I(_01369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05847__A1 (.I(_01369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05833__A1 (.I(_01369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04882__I (.I(_01369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04857__A1 (.I(_01369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04845__A1 (.I(_01369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07738__C (.I(_01370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06484__A2 (.I(_01370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05892__A1 (.I(_01370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05885__A2 (.I(_01370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05882__A2 (.I(_01370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05872__A1 (.I(_01370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05852__A1 (.I(_01370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05849__I (.I(_01370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04883__A1 (.I(_01370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04857__A2 (.I(_01370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04845__A2 (.I(_01370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08625__A1 (.I(_01372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08424__A1 (.I(_01372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08219__A1 (.I(_01372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06476__A1 (.I(_01372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05979__A1 (.I(_01372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05967__A1 (.I(_01372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05910__A1 (.I(_01372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05883__B (.I(_01372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05833__A2 (.I(_01372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05830__A1 (.I(_01372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04852__A1 (.I(_01372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04847__I (.I(_01372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08445__A1 (.I(_01373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06486__A1 (.I(_01373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05992__C (.I(_01373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05908__A1 (.I(_01373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05893__B (.I(_01373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05885__A1 (.I(_01373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04850__A1 (.I(_01373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08515__A1 (.I(_01374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08228__A1 (.I(_01374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07741__C (.I(_01374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05973__A1 (.I(_01374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05972__A1 (.I(_01374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05967__A2 (.I(_01374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05929__A1 (.I(_01374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05928__A1 (.I(_01374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05926__A1 (.I(_01374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05920__A1 (.I(_01374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05915__A1 (.I(_01374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05900__A1 (.I(_01374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05833__A3 (.I(_01374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05824__C (.I(_01374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04852__A2 (.I(_01374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04849__I (.I(_01374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09373__C (.I(_01375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09369__A1 (.I(_01375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08513__A1 (.I(_01375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06486__C (.I(_01375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05976__A1 (.I(_01375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05880__A4 (.I(_01375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04850__A2 (.I(_01375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09391__A2 (.I(_01377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04887__C (.I(_01377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04878__A1 (.I(_01377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04862__A2 (.I(_01377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09377__A1 (.I(_01381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08264__A1 (.I(_01381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05920__B1 (.I(_01381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04856__B (.I(_01381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09369__B2 (.I(_01385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09365__A1 (.I(_01385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06487__A2 (.I(_01385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05880__A3 (.I(_01385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04860__C (.I(_01385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09380__B (.I(_01386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09360__A2 (.I(_01386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08723__A2 (.I(_01386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06230__A1 (.I(_01386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06159__A2 (.I(_01386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06006__A1 (.I(_01386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06000__A2 (.I(_01386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05999__A1 (.I(_01386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05930__A1 (.I(_01386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05929__C (.I(_01386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05867__A2 (.I(_01386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04861__B (.I(_01386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05990__A1 (.I(_01387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04888__A2 (.I(_01387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04878__A2 (.I(_01387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04869__B (.I(_01387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04862__A3 (.I(_01387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04898__A2 (.I(_01388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04894__A2 (.I(_01388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04875__A2 (.I(_01388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04863__A2 (.I(_01388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08473__A1 (.I(_01390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05847__A2 (.I(_01390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04865__A1 (.I(_01390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09391__B (.I(_01393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09373__A2 (.I(_01393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05994__A1 (.I(_01393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05866__A1 (.I(_01393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04869__A1 (.I(_01393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05999__A2 (.I(_01394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04869__A2 (.I(_01394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05762__A1 (.I(_01397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05674__A1 (.I(_01397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05586__A1 (.I(_01397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05498__A1 (.I(_01397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05144__I (.I(_01397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05122__I (.I(_01397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05105__I (.I(_01397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05097__I (.I(_01397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05061__I (.I(_01397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04872__I (.I(_01397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05790__A1 (.I(_01398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05735__A1 (.I(_01398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05702__A1 (.I(_01398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05614__A1 (.I(_01398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05526__A1 (.I(_01398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05516__A1 (.I(_01398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05438__A1 (.I(_01398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05428__A1 (.I(_01398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05350__A1 (.I(_01398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05340__A1 (.I(_01398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05262__A1 (.I(_01398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05252__A1 (.I(_01398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05167__A1 (.I(_01398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05152__A1 (.I(_01398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05078__I (.I(_01398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04873__I (.I(_01398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05810__A1 (.I(_01399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05726__A1 (.I(_01399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05722__A1 (.I(_01399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05638__A1 (.I(_01399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05634__A1 (.I(_01399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05550__A1 (.I(_01399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05546__A1 (.I(_01399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05462__A1 (.I(_01399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05458__A1 (.I(_01399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05374__A1 (.I(_01399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05370__A1 (.I(_01399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05286__A1 (.I(_01399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05282__A1 (.I(_01399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05198__A1 (.I(_01399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05191__A1 (.I(_01399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04902__A1 (.I(_01399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05808__B (.I(_01402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05720__B (.I(_01402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05632__B (.I(_01402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05544__B (.I(_01402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05456__B (.I(_01402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05368__B (.I(_01402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05280__B (.I(_01402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05187__B (.I(_01402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04879__A1 (.I(_01402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05963__A1 (.I(_01403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05962__A2 (.I(_01403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05961__A1 (.I(_01403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05960__A2 (.I(_01403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05959__A1 (.I(_01403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05958__A2 (.I(_01403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05957__A1 (.I(_01403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05956__A2 (.I(_01403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05955__A1 (.I(_01403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05954__A2 (.I(_01403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05953__A1 (.I(_01403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05952__A2 (.I(_01403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05951__A1 (.I(_01403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05950__A2 (.I(_01403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04903__I (.I(_01403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04878__B (.I(_01403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05817__C (.I(_01404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05729__C (.I(_01404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05641__C (.I(_01404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05553__C (.I(_01404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05465__C (.I(_01404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05377__C (.I(_01404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05289__C (.I(_01404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05201__C (.I(_01404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04879__A2 (.I(_01404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05819__A1 (.I(_01406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05731__A1 (.I(_01406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05643__A1 (.I(_01406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05555__A1 (.I(_01406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05467__A1 (.I(_01406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05379__A1 (.I(_01406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05291__A1 (.I(_01406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05203__A1 (.I(_01406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04901__A1 (.I(_01406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08253__A1 (.I(_01408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07737__A1 (.I(_01408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06484__A1 (.I(_01408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04884__A1 (.I(_01408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05965__B1 (.I(_01409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05903__B2 (.I(_01409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05883__A1 (.I(_01409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05865__A1 (.I(_01409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05823__I (.I(_01409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04884__A2 (.I(_01409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08722__A2 (.I(_01410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05878__A1 (.I(_01410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04885__A1 (.I(_01410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05861__A3 (.I(_01411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05856__A2 (.I(_01411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04887__A1 (.I(_01411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06005__A2 (.I(_01412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04887__A2 (.I(_01412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05072__A2 (.I(_01414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04889__A2 (.I(_01414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05773__B (.I(_01416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05762__B (.I(_01416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05685__B (.I(_01416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05674__B (.I(_01416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05597__B (.I(_01416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05509__B (.I(_01416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05421__B (.I(_01416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05333__B (.I(_01416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05245__B (.I(_01416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05156__I (.I(_01416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05143__B (.I(_01416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05113__I (.I(_01416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04891__I (.I(_01416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05748__B (.I(_01417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05735__B (.I(_01417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05647__B (.I(_01417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05629__B (.I(_01417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05559__B (.I(_01417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05541__B (.I(_01417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05471__B (.I(_01417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05453__B (.I(_01417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05383__B (.I(_01417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05365__B (.I(_01417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05295__B (.I(_01417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05277__B (.I(_01417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05207__B (.I(_01417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05184__B (.I(_01417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05067__B (.I(_01417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04892__I (.I(_01417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05816__B (.I(_01418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05728__B (.I(_01418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05660__B (.I(_01418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05640__B (.I(_01418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05572__B (.I(_01418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05552__B (.I(_01418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05484__B (.I(_01418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05464__B (.I(_01418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05396__B (.I(_01418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05376__B (.I(_01418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05308__B (.I(_01418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05288__B (.I(_01418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05220__B (.I(_01418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05200__B (.I(_01418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05095__B (.I(_01418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04901__A2 (.I(_01418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05047__A1 (.I(_01419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04895__A1 (.I(_01419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05047__A2 (.I(_01420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04895__A2 (.I(_01420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05768__A1 (.I(_01421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04896__I (.I(_01421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05788__A1 (.I(_01422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05700__A1 (.I(_01422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05680__A1 (.I(_01422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05612__A1 (.I(_01422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05592__A1 (.I(_01422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05524__A1 (.I(_01422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05504__A1 (.I(_01422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05436__A1 (.I(_01422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05416__A1 (.I(_01422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05348__A1 (.I(_01422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05328__A1 (.I(_01422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05260__A1 (.I(_01422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05240__A1 (.I(_01422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05165__A1 (.I(_01422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05138__A1 (.I(_01422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04901__A3 (.I(_01422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05758__C (.I(_01425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05115__I (.I(_01425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04900__I (.I(_01425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05749__C (.I(_01426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05709__C (.I(_01426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05661__C (.I(_01426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05621__C (.I(_01426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05573__C (.I(_01426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05533__C (.I(_01426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05485__C (.I(_01426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05445__C (.I(_01426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05397__C (.I(_01426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05357__C (.I(_01426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05309__C (.I(_01426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05269__C (.I(_01426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05221__C (.I(_01426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05174__C (.I(_01426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05096__C (.I(_01426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04901__A4 (.I(_01426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09398__A1 (.I(_01428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08923__A1 (.I(_01428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08656__A1 (.I(_01428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08654__B (.I(_01428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07746__A1 (.I(_01428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07730__A1 (.I(_01428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07689__A1 (.I(_01428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07682__A1 (.I(_01428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07681__A1 (.I(_01428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07676__A1 (.I(_01428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07672__A1 (.I(_01428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06473__A1 (.I(_01428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04905__I (.I(_01428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09567__A1 (.I(_01429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09388__B (.I(_01429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07690__A1 (.I(_01429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07687__A1 (.I(_01429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07685__C (.I(_01429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07677__B (.I(_01429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04919__A1 (.I(_01429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04906__A1 (.I(_01429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08197__A2 (.I(_01431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06469__A2 (.I(_01431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05971__A2 (.I(_01431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05045__S (.I(_01431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04938__A1 (.I(_01431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04918__A1 (.I(_01431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04910__A2 (.I(_01431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04908__A2 (.I(_01431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08144__S (.I(_01434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08142__S (.I(_01434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08141__S (.I(_01434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04932__A1 (.I(_01434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04913__I (.I(_01434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08235__S (.I(_01435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08188__S (.I(_01435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08184__A1 (.I(_01435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08177__A1 (.I(_01435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08175__S (.I(_01435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08172__S (.I(_01435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08166__A1 (.I(_01435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08163__S (.I(_01435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08162__S (.I(_01435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08161__A1 (.I(_01435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08160__A1 (.I(_01435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08156__S (.I(_01435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08155__S (.I(_01435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08143__S (.I(_01435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06468__I (.I(_01435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04914__I (.I(_01435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08488__S (.I(_01436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08474__S (.I(_01436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08429__A1 (.I(_01436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08400__A1 (.I(_01436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08346__S (.I(_01436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08309__S (.I(_01436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08307__S (.I(_01436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08277__S (.I(_01436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08203__S (.I(_01436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08200__A1 (.I(_01436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08168__S (.I(_01436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08158__A1 (.I(_01436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08153__A1 (.I(_01436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08150__A1 (.I(_01436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08146__A1 (.I(_01436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04915__I (.I(_01436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08922__A1 (.I(_01437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08519__S (.I(_01437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08510__A1 (.I(_01437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08509__A1 (.I(_01437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08498__S (.I(_01437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08415__S (.I(_01437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08407__A1 (.I(_01437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08395__A1 (.I(_01437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08390__S (.I(_01437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08376__A1 (.I(_01437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08359__S (.I(_01437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08265__S (.I(_01437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08254__S (.I(_01437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04928__A1 (.I(_01437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04917__A1 (.I(_01437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04916__A1 (.I(_01437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08012__A2 (.I(_01442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06485__A2 (.I(_01442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05013__A2 (.I(_01442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05008__A2 (.I(_01442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04995__A2 (.I(_01442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04991__A2 (.I(_01442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04984__A2 (.I(_01442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04980__A2 (.I(_01442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04974__B (.I(_01442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04971__A2 (.I(_01442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04958__B (.I(_01442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04939__I (.I(_01442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04924__I (.I(_01442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04921__I (.I(_01442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05041__A1 (.I(_01443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05037__A1 (.I(_01443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05014__A1 (.I(_01443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05009__A1 (.I(_01443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04996__A1 (.I(_01443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04992__A1 (.I(_01443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04985__A1 (.I(_01443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04981__A1 (.I(_01443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04973__A2 (.I(_01443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04972__A1 (.I(_01443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04965__A1 (.I(_01443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04955__A2 (.I(_01443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04934__A2 (.I(_01443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04930__A2 (.I(_01443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04926__A2 (.I(_01443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04922__A2 (.I(_01443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05969__B (.I(_01445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05033__A1 (.I(_01445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05029__A1 (.I(_01445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05025__A1 (.I(_01445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05021__A1 (.I(_01445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05017__A1 (.I(_01445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05003__A1 (.I(_01445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04999__A1 (.I(_01445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04988__A1 (.I(_01445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04968__A1 (.I(_01445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04954__A1 (.I(_01445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04951__A1 (.I(_01445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04944__A1 (.I(_01445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04935__A1 (.I(_01445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04931__A1 (.I(_01445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04927__A1 (.I(_01445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05040__A2 (.I(_01457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05036__A2 (.I(_01457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05032__A2 (.I(_01457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05028__A2 (.I(_01457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05024__A2 (.I(_01457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05020__A2 (.I(_01457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05016__A2 (.I(_01457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05002__A2 (.I(_01457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04998__A2 (.I(_01457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04987__A2 (.I(_01457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04967__A2 (.I(_01457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04964__A2 (.I(_01457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04953__A2 (.I(_01457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04950__A2 (.I(_01457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04943__A2 (.I(_01457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04940__A2 (.I(_01457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04963__A3 (.I(_01462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04948__A2 (.I(_01462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04947__A2 (.I(_01462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05046__I (.I(_01538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05807__A1 (.I(_01539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05769__A1 (.I(_01539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05719__A1 (.I(_01539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05681__A1 (.I(_01539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05631__A1 (.I(_01539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05593__A1 (.I(_01539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05543__A1 (.I(_01539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05505__A1 (.I(_01539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05455__A1 (.I(_01539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05417__A1 (.I(_01539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05367__A1 (.I(_01539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05329__A1 (.I(_01539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05279__A1 (.I(_01539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05241__A1 (.I(_01539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05186__A1 (.I(_01539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05139__A1 (.I(_01539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05753__A1 (.I(_01540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05665__A1 (.I(_01540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05577__A1 (.I(_01540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05175__I (.I(_01540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05153__I (.I(_01540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05117__I (.I(_01540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05109__I (.I(_01540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05102__I (.I(_01540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05049__I (.I(_01540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05794__A1 (.I(_01541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05784__A1 (.I(_01541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05696__A1 (.I(_01541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05608__A1 (.I(_01541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05520__A1 (.I(_01541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05502__A1 (.I(_01541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05432__A1 (.I(_01541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05414__A1 (.I(_01541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05344__A1 (.I(_01541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05326__A1 (.I(_01541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05256__A1 (.I(_01541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05238__A1 (.I(_01541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05159__A1 (.I(_01541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05135__A1 (.I(_01541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05070__I (.I(_01541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05050__I (.I(_01541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05748__A1 (.I(_01542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05733__A1 (.I(_01542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05660__A1 (.I(_01542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05645__A1 (.I(_01542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05572__A1 (.I(_01542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05557__A1 (.I(_01542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05484__A1 (.I(_01542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05469__A1 (.I(_01542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05396__A1 (.I(_01542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05381__A1 (.I(_01542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05308__A1 (.I(_01542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05293__A1 (.I(_01542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05220__A1 (.I(_01542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05205__A1 (.I(_01542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05095__A1 (.I(_01542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05060__A1 (.I(_01542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06070__B (.I(_01543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06009__A1 (.I(_01543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05123__I (.I(_01543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05110__I (.I(_01543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05085__I (.I(_01543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05063__I (.I(_01543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05052__I (.I(_01543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05752__S0 (.I(_01544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05664__S0 (.I(_01544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05576__S0 (.I(_01544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05488__S0 (.I(_01544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05400__S0 (.I(_01544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05312__S0 (.I(_01544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05224__S0 (.I(_01544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05154__I (.I(_01544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05131__I (.I(_01544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05127__I (.I(_01544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05118__I (.I(_01544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05106__I (.I(_01544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05103__S0 (.I(_01544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05098__I (.I(_01544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05079__I (.I(_01544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05053__I (.I(_01544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05779__S0 (.I(_01545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05759__S0 (.I(_01545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05691__S0 (.I(_01545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05671__S0 (.I(_01545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05603__S0 (.I(_01545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05583__S0 (.I(_01545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05515__S0 (.I(_01545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05495__S0 (.I(_01545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05427__S0 (.I(_01545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05407__S0 (.I(_01545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05339__S0 (.I(_01545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05265__S0 (.I(_01545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05251__S0 (.I(_01545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05170__S0 (.I(_01545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05151__S0 (.I(_01545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05054__I (.I(_01545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05745__S0 (.I(_01546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05732__S0 (.I(_01546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05657__S0 (.I(_01546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05644__S0 (.I(_01546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05560__S0 (.I(_01546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05556__S0 (.I(_01546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05472__S0 (.I(_01546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05468__S0 (.I(_01546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05384__S0 (.I(_01546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05380__S0 (.I(_01546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05296__S0 (.I(_01546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05292__S0 (.I(_01546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05208__S0 (.I(_01546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05204__S0 (.I(_01546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05068__S0 (.I(_01546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05059__S0 (.I(_01546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06071__A1 (.I(_01547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05160__I (.I(_01547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05132__I (.I(_01547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05124__I (.I(_01547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05111__I (.I(_01547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05087__I (.I(_01547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05056__I (.I(_01547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05752__S1 (.I(_01548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05664__S1 (.I(_01548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05576__S1 (.I(_01548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05488__S1 (.I(_01548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05400__S1 (.I(_01548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05312__S1 (.I(_01548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05224__S1 (.I(_01548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05176__I (.I(_01548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05150__I (.I(_01548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05128__I (.I(_01548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05119__I (.I(_01548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05103__S1 (.I(_01548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05099__I (.I(_01548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05081__I (.I(_01548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05065__I (.I(_01548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05057__I (.I(_01548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05804__S1 (.I(_01549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05774__S1 (.I(_01549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05716__S1 (.I(_01549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05686__S1 (.I(_01549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05628__S1 (.I(_01549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05598__S1 (.I(_01549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05540__S1 (.I(_01549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05510__S1 (.I(_01549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05452__S1 (.I(_01549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05422__S1 (.I(_01549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05364__S1 (.I(_01549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05334__S1 (.I(_01549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05276__S1 (.I(_01549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05183__S1 (.I(_01549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05179__S1 (.I(_01549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05058__I (.I(_01549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05745__S1 (.I(_01550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05732__S1 (.I(_01550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05648__S1 (.I(_01550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05644__S1 (.I(_01550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05560__S1 (.I(_01550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05556__S1 (.I(_01550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05472__S1 (.I(_01550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05468__S1 (.I(_01550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05384__S1 (.I(_01550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05380__S1 (.I(_01550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05296__S1 (.I(_01550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05292__S1 (.I(_01550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05208__S1 (.I(_01550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05204__S1 (.I(_01550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05068__S1 (.I(_01550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05059__S1 (.I(_01550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05060__A2 (.I(_01551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05805__A1 (.I(_01553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05801__A1 (.I(_01553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05717__A1 (.I(_01553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05713__A1 (.I(_01553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05629__A1 (.I(_01553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05625__A1 (.I(_01553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05537__A1 (.I(_01553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05449__A1 (.I(_01553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05444__A1 (.I(_01553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05361__A1 (.I(_01553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05356__A1 (.I(_01553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05273__A1 (.I(_01553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05268__A1 (.I(_01553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05180__A1 (.I(_01553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05173__A1 (.I(_01553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05062__I (.I(_01553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05746__A1 (.I(_01554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05737__A1 (.I(_01554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05649__A1 (.I(_01554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05647__A1 (.I(_01554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05561__A1 (.I(_01554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05559__A1 (.I(_01554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05473__A1 (.I(_01554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05471__A1 (.I(_01554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05385__A1 (.I(_01554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05383__A1 (.I(_01554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05297__A1 (.I(_01554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05295__A1 (.I(_01554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05209__A1 (.I(_01554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05207__A1 (.I(_01554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05069__A1 (.I(_01554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05067__A1 (.I(_01554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05800__S0 (.I(_01555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05795__S0 (.I(_01555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05712__S0 (.I(_01555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05707__S0 (.I(_01555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05624__S0 (.I(_01555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05619__S0 (.I(_01555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05536__S0 (.I(_01555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05531__S0 (.I(_01555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05448__S0 (.I(_01555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05443__S0 (.I(_01555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05360__S0 (.I(_01555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05355__S0 (.I(_01555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05272__S0 (.I(_01555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05267__S0 (.I(_01555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05172__S0 (.I(_01555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05064__I (.I(_01555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05743__S0 (.I(_01556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05738__S0 (.I(_01556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05655__S0 (.I(_01556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05650__S0 (.I(_01556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05562__S0 (.I(_01556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05558__S0 (.I(_01556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05474__S0 (.I(_01556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05470__S0 (.I(_01556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05386__S0 (.I(_01556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05382__S0 (.I(_01556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05298__S0 (.I(_01556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05294__S0 (.I(_01556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05210__S0 (.I(_01556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05206__S0 (.I(_01556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05071__S0 (.I(_01556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05066__S0 (.I(_01556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05743__S1 (.I(_01557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05738__S1 (.I(_01557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05650__S1 (.I(_01557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05646__S1 (.I(_01557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05562__S1 (.I(_01557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05558__S1 (.I(_01557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05474__S1 (.I(_01557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05470__S1 (.I(_01557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05386__S1 (.I(_01557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05382__S1 (.I(_01557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05298__S1 (.I(_01557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05294__S1 (.I(_01557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05210__S1 (.I(_01557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05206__S1 (.I(_01557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05071__S1 (.I(_01557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05066__S1 (.I(_01557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05069__A2 (.I(_01560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05744__A1 (.I(_01562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05739__A1 (.I(_01562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05656__A1 (.I(_01562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05651__A1 (.I(_01562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05568__A1 (.I(_01562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05563__A1 (.I(_01562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05480__A1 (.I(_01562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05475__A1 (.I(_01562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05392__A1 (.I(_01562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05387__A1 (.I(_01562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05304__A1 (.I(_01562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05299__A1 (.I(_01562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05216__A1 (.I(_01562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05211__A1 (.I(_01562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05091__A1 (.I(_01562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05074__A1 (.I(_01562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05777__B (.I(_01564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05753__B (.I(_01564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05665__B (.I(_01564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05577__B (.I(_01564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05489__B (.I(_01564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05401__B (.I(_01564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05313__B (.I(_01564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05225__B (.I(_01564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05162__I (.I(_01564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05134__I (.I(_01564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05104__B (.I(_01564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05073__I (.I(_01564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05739__B (.I(_01565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05713__B (.I(_01565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05651__B (.I(_01565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05625__B (.I(_01565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05563__B (.I(_01565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05537__B (.I(_01565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05475__B (.I(_01565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05449__B (.I(_01565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05387__B (.I(_01565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05361__B (.I(_01565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05299__B (.I(_01565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05273__B (.I(_01565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05211__B (.I(_01565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05180__B (.I(_01565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05090__I (.I(_01565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05074__B (.I(_01565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05136__I (.I(_01567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05076__I (.I(_01567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05806__C (.I(_01568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05740__C (.I(_01568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05718__C (.I(_01568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05652__C (.I(_01568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05630__C (.I(_01568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05564__C (.I(_01568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05542__C (.I(_01568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05476__C (.I(_01568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05454__C (.I(_01568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05388__C (.I(_01568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05366__C (.I(_01568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05300__C (.I(_01568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05278__C (.I(_01568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05212__C (.I(_01568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05185__C (.I(_01568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05077__C (.I(_01568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05139__A2 (.I(_01569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05814__A1 (.I(_01570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05742__A1 (.I(_01570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05658__A1 (.I(_01570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05654__A1 (.I(_01570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05570__A1 (.I(_01570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05566__A1 (.I(_01570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05482__A1 (.I(_01570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05478__A1 (.I(_01570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05394__A1 (.I(_01570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05390__A1 (.I(_01570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05306__A1 (.I(_01570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05302__A1 (.I(_01570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05218__A1 (.I(_01570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05214__A1 (.I(_01570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05093__A1 (.I(_01570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05084__A1 (.I(_01570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05798__S0 (.I(_01571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05734__S0 (.I(_01571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05710__S0 (.I(_01571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05646__S0 (.I(_01571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05622__S0 (.I(_01571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05534__S0 (.I(_01571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05446__S0 (.I(_01571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05362__S0 (.I(_01571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05358__S0 (.I(_01571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05274__S0 (.I(_01571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05270__S0 (.I(_01571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05195__I (.I(_01571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05188__I (.I(_01571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05181__S0 (.I(_01571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05177__S0 (.I(_01571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05080__I (.I(_01571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05813__S0 (.I(_01572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05741__S0 (.I(_01572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05725__S0 (.I(_01572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05653__S0 (.I(_01572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05569__S0 (.I(_01572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05565__S0 (.I(_01572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05481__S0 (.I(_01572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05477__S0 (.I(_01572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05393__S0 (.I(_01572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05389__S0 (.I(_01572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05305__S0 (.I(_01572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05301__S0 (.I(_01572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05217__S0 (.I(_01572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05213__S0 (.I(_01572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05092__S0 (.I(_01572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05083__S0 (.I(_01572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05770__S1 (.I(_01573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05754__S1 (.I(_01573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05682__S1 (.I(_01573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05666__S1 (.I(_01573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05594__S1 (.I(_01573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05578__S1 (.I(_01573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05506__S1 (.I(_01573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05490__S1 (.I(_01573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05418__S1 (.I(_01573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05402__S1 (.I(_01573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05314__S1 (.I(_01573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05246__S1 (.I(_01573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05226__S1 (.I(_01573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05145__S1 (.I(_01573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05107__S1 (.I(_01573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05082__I (.I(_01573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05813__S1 (.I(_01574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05741__S1 (.I(_01574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05657__S1 (.I(_01574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05653__S1 (.I(_01574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05569__S1 (.I(_01574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05565__S1 (.I(_01574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05481__S1 (.I(_01574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05477__S1 (.I(_01574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05393__S1 (.I(_01574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05389__S1 (.I(_01574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05305__S1 (.I(_01574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05301__S1 (.I(_01574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05217__S1 (.I(_01574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05213__S1 (.I(_01574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05092__S1 (.I(_01574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05083__S1 (.I(_01574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05084__A2 (.I(_01575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05804__S0 (.I(_01577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05774__S0 (.I(_01577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05716__S0 (.I(_01577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05686__S0 (.I(_01577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05628__S0 (.I(_01577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05598__S0 (.I(_01577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05540__S0 (.I(_01577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05510__S0 (.I(_01577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05452__S0 (.I(_01577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05422__S0 (.I(_01577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05364__S0 (.I(_01577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05334__S0 (.I(_01577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05276__S0 (.I(_01577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05183__S0 (.I(_01577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05179__S0 (.I(_01577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05086__I (.I(_01577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05747__S0 (.I(_01578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05736__S0 (.I(_01578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05659__S0 (.I(_01578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05648__S0 (.I(_01578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05571__S0 (.I(_01578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05567__S0 (.I(_01578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05483__S0 (.I(_01578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05479__S0 (.I(_01578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05395__S0 (.I(_01578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05391__S0 (.I(_01578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05307__S0 (.I(_01578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05303__S0 (.I(_01578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05219__S0 (.I(_01578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05215__S0 (.I(_01578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05094__S0 (.I(_01578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05089__S0 (.I(_01578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05776__S1 (.I(_01579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05756__S1 (.I(_01579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05688__S1 (.I(_01579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05668__S1 (.I(_01579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05600__S1 (.I(_01579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05580__S1 (.I(_01579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05512__S1 (.I(_01579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05492__S1 (.I(_01579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05424__S1 (.I(_01579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05404__S1 (.I(_01579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05336__S1 (.I(_01579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05316__S1 (.I(_01579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05248__S1 (.I(_01579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05228__S1 (.I(_01579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05147__S1 (.I(_01579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05088__I (.I(_01579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05747__S1 (.I(_01580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05736__S1 (.I(_01580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05659__S1 (.I(_01580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05655__S1 (.I(_01580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05571__S1 (.I(_01580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05567__S1 (.I(_01580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05483__S1 (.I(_01580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05479__S1 (.I(_01580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05395__S1 (.I(_01580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05391__S1 (.I(_01580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05307__S1 (.I(_01580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05303__S1 (.I(_01580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05219__S1 (.I(_01580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05215__S1 (.I(_01580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05094__S1 (.I(_01580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05089__S1 (.I(_01580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05091__A2 (.I(_01581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05812__B (.I(_01582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05744__B (.I(_01582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05724__B (.I(_01582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05656__B (.I(_01582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05636__B (.I(_01582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05568__B (.I(_01582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05548__B (.I(_01582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05480__B (.I(_01582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05460__B (.I(_01582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05392__B (.I(_01582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05372__B (.I(_01582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05304__B (.I(_01582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05284__B (.I(_01582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05216__B (.I(_01582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05194__B (.I(_01582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05091__B (.I(_01582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05093__A2 (.I(_01584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05095__A2 (.I(_01586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05139__A3 (.I(_01588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05780__A1 (.I(_01589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05751__A1 (.I(_01589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05692__A1 (.I(_01589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05663__A1 (.I(_01589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05604__A1 (.I(_01589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05575__A1 (.I(_01589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05500__A1 (.I(_01589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05487__A1 (.I(_01589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05412__A1 (.I(_01589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05399__A1 (.I(_01589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05324__A1 (.I(_01589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05311__A1 (.I(_01589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05236__A1 (.I(_01589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05223__A1 (.I(_01589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05130__A1 (.I(_01589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05101__A1 (.I(_01589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05793__S0 (.I(_01590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05750__S0 (.I(_01590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05705__S0 (.I(_01590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05662__S0 (.I(_01590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05617__S0 (.I(_01590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05574__S0 (.I(_01590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05529__S0 (.I(_01590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05486__S0 (.I(_01590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05441__S0 (.I(_01590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05398__S0 (.I(_01590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05353__S0 (.I(_01590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05310__S0 (.I(_01590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05255__S0 (.I(_01590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05222__S0 (.I(_01590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05158__S0 (.I(_01590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05100__S0 (.I(_01590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06011__A1 (.I(_01591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05793__S1 (.I(_01591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05750__S1 (.I(_01591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05705__S1 (.I(_01591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05662__S1 (.I(_01591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05617__S1 (.I(_01591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05574__S1 (.I(_01591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05529__S1 (.I(_01591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05486__S1 (.I(_01591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05398__S1 (.I(_01591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05343__S1 (.I(_01591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05310__S1 (.I(_01591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05255__S1 (.I(_01591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05222__S1 (.I(_01591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05158__S1 (.I(_01591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05100__S1 (.I(_01591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05116__A1 (.I(_01593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05777__A1 (.I(_01594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05773__A1 (.I(_01594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05689__A1 (.I(_01594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05685__A1 (.I(_01594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05601__A1 (.I(_01594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05597__A1 (.I(_01594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05509__A1 (.I(_01594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05489__A1 (.I(_01594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05421__A1 (.I(_01594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05401__A1 (.I(_01594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05333__A1 (.I(_01594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05313__A1 (.I(_01594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05245__A1 (.I(_01594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05225__A1 (.I(_01594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05143__A1 (.I(_01594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05104__A1 (.I(_01594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05104__A2 (.I(_01595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05771__A1 (.I(_01597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05764__A1 (.I(_01597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05683__A1 (.I(_01597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05676__A1 (.I(_01597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05595__A1 (.I(_01597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05588__A1 (.I(_01597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05507__A1 (.I(_01597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05491__A1 (.I(_01597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05419__A1 (.I(_01597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05403__A1 (.I(_01597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05331__A1 (.I(_01597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05315__A1 (.I(_01597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05243__A1 (.I(_01597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05227__A1 (.I(_01597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05141__A1 (.I(_01597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05108__A1 (.I(_01597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05770__S0 (.I(_01598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05754__S0 (.I(_01598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05682__S0 (.I(_01598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05666__S0 (.I(_01598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05594__S0 (.I(_01598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05578__S0 (.I(_01598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05506__S0 (.I(_01598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05490__S0 (.I(_01598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05418__S0 (.I(_01598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05402__S0 (.I(_01598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05330__S0 (.I(_01598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05314__S0 (.I(_01598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05246__S0 (.I(_01598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05226__S0 (.I(_01598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05145__S0 (.I(_01598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05107__S0 (.I(_01598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05108__A2 (.I(_01599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05782__A1 (.I(_01601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05757__A1 (.I(_01601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05694__A1 (.I(_01601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05669__A1 (.I(_01601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05606__A1 (.I(_01601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05581__A1 (.I(_01601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05513__A1 (.I(_01601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05493__A1 (.I(_01601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05425__A1 (.I(_01601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05405__A1 (.I(_01601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05337__A1 (.I(_01601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05317__A1 (.I(_01601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05249__A1 (.I(_01601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05229__A1 (.I(_01601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05148__A1 (.I(_01601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05114__A1 (.I(_01601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05776__S0 (.I(_01602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05756__S0 (.I(_01602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05688__S0 (.I(_01602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05668__S0 (.I(_01602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05600__S0 (.I(_01602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05580__S0 (.I(_01602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05512__S0 (.I(_01602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05492__S0 (.I(_01602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05424__S0 (.I(_01602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05404__S0 (.I(_01602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05336__S0 (.I(_01602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05316__S0 (.I(_01602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05248__S0 (.I(_01602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05228__S0 (.I(_01602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05147__S0 (.I(_01602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05112__S0 (.I(_01602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05791__S1 (.I(_01603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05781__S1 (.I(_01603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05703__S1 (.I(_01603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05693__S1 (.I(_01603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05615__S1 (.I(_01603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05605__S1 (.I(_01603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05527__S1 (.I(_01603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05517__S1 (.I(_01603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05439__S1 (.I(_01603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05429__S1 (.I(_01603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05351__S1 (.I(_01603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05341__S1 (.I(_01603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05263__S1 (.I(_01603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05253__S1 (.I(_01603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05155__S1 (.I(_01603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05112__S1 (.I(_01603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05114__A2 (.I(_01604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05782__B (.I(_01605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05757__B (.I(_01605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05694__B (.I(_01605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05669__B (.I(_01605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05586__B (.I(_01605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05581__B (.I(_01605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05498__B (.I(_01605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05493__B (.I(_01605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05410__B (.I(_01605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05405__B (.I(_01605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05322__B (.I(_01605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05317__B (.I(_01605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05234__B (.I(_01605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05229__B (.I(_01605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05126__B (.I(_01605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05114__B (.I(_01605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05797__C (.I(_01607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05787__C (.I(_01607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05699__C (.I(_01607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05670__C (.I(_01607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05611__C (.I(_01607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05582__C (.I(_01607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05523__C (.I(_01607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05494__C (.I(_01607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05435__C (.I(_01607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05406__C (.I(_01607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05347__C (.I(_01607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05318__C (.I(_01607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05259__C (.I(_01607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05230__C (.I(_01607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05164__C (.I(_01607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05116__C (.I(_01607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05803__A1 (.I(_01609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05760__A1 (.I(_01609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05706__A1 (.I(_01609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05672__A1 (.I(_01609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05618__A1 (.I(_01609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05584__A1 (.I(_01609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05530__A1 (.I(_01609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05496__A1 (.I(_01609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05442__A1 (.I(_01609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05408__A1 (.I(_01609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05354__A1 (.I(_01609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05320__A1 (.I(_01609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05266__A1 (.I(_01609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05232__A1 (.I(_01609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05171__A1 (.I(_01609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05121__A1 (.I(_01609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05802__S0 (.I(_01610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05789__S0 (.I(_01610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05714__S0 (.I(_01610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05701__S0 (.I(_01610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05626__S0 (.I(_01610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05613__S0 (.I(_01610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05538__S0 (.I(_01610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05525__S0 (.I(_01610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05450__S0 (.I(_01610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05437__S0 (.I(_01610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05349__S0 (.I(_01610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05319__S0 (.I(_01610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05261__S0 (.I(_01610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05231__S0 (.I(_01610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05166__S0 (.I(_01610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05120__S0 (.I(_01610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05802__S1 (.I(_01611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05789__S1 (.I(_01611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05714__S1 (.I(_01611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05701__S1 (.I(_01611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05626__S1 (.I(_01611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05613__S1 (.I(_01611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05538__S1 (.I(_01611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05525__S1 (.I(_01611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05437__S1 (.I(_01611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05407__S1 (.I(_01611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05349__S1 (.I(_01611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05319__S1 (.I(_01611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05261__S1 (.I(_01611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05231__S1 (.I(_01611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05166__S1 (.I(_01611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05120__S1 (.I(_01611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05121__A2 (.I(_01612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05796__A1 (.I(_01614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05786__A1 (.I(_01614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05708__A1 (.I(_01614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05698__A1 (.I(_01614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05620__A1 (.I(_01614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05610__A1 (.I(_01614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05532__A1 (.I(_01614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05522__A1 (.I(_01614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05434__A1 (.I(_01614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05410__A1 (.I(_01614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05346__A1 (.I(_01614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05322__A1 (.I(_01614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05258__A1 (.I(_01614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05234__A1 (.I(_01614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05163__A1 (.I(_01614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05126__A1 (.I(_01614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05772__S0 (.I(_01615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05761__S0 (.I(_01615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05684__S0 (.I(_01615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05673__S0 (.I(_01615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05596__S0 (.I(_01615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05585__S0 (.I(_01615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05508__S0 (.I(_01615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05497__S0 (.I(_01615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05420__S0 (.I(_01615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05409__S0 (.I(_01615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05332__S0 (.I(_01615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05321__S0 (.I(_01615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05244__S0 (.I(_01615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05233__S0 (.I(_01615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05142__S0 (.I(_01615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05125__S0 (.I(_01615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05772__S1 (.I(_01616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05761__S1 (.I(_01616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05684__S1 (.I(_01616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05673__S1 (.I(_01616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05596__S1 (.I(_01616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05585__S1 (.I(_01616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05508__S1 (.I(_01616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05497__S1 (.I(_01616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05420__S1 (.I(_01616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05409__S1 (.I(_01616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05332__S1 (.I(_01616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05321__S1 (.I(_01616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05244__S1 (.I(_01616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05233__S1 (.I(_01616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05142__S1 (.I(_01616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05125__S1 (.I(_01616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05126__A2 (.I(_01617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05137__A2 (.I(_01618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05783__S0 (.I(_01619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05763__S0 (.I(_01619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05695__S0 (.I(_01619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05675__S0 (.I(_01619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05607__S0 (.I(_01619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05587__S0 (.I(_01619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05519__S0 (.I(_01619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05499__S0 (.I(_01619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05431__S0 (.I(_01619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05411__S0 (.I(_01619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05343__S0 (.I(_01619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05323__S0 (.I(_01619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05242__S0 (.I(_01619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05235__S0 (.I(_01619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05140__S0 (.I(_01619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05129__S0 (.I(_01619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05783__S1 (.I(_01620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05763__S1 (.I(_01620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05695__S1 (.I(_01620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05675__S1 (.I(_01620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05607__S1 (.I(_01620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05587__S1 (.I(_01620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05519__S1 (.I(_01620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05499__S1 (.I(_01620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05431__S1 (.I(_01620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05411__S1 (.I(_01620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05330__S1 (.I(_01620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05323__S1 (.I(_01620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05242__S1 (.I(_01620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05235__S1 (.I(_01620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05140__S1 (.I(_01620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05129__S1 (.I(_01620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05785__S0 (.I(_01623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05765__S0 (.I(_01623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05697__S0 (.I(_01623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05677__S0 (.I(_01623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05609__S0 (.I(_01623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05589__S0 (.I(_01623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05521__S0 (.I(_01623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05501__S0 (.I(_01623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05433__S0 (.I(_01623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05413__S0 (.I(_01623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05345__S0 (.I(_01623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05325__S0 (.I(_01623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05257__S0 (.I(_01623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05237__S0 (.I(_01623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05161__S0 (.I(_01623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05133__S0 (.I(_01623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05785__S1 (.I(_01624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05765__S1 (.I(_01624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05697__S1 (.I(_01624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05677__S1 (.I(_01624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05609__S1 (.I(_01624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05589__S1 (.I(_01624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05521__S1 (.I(_01624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05501__S1 (.I(_01624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05433__S1 (.I(_01624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05413__S1 (.I(_01624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05345__S1 (.I(_01624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05325__S1 (.I(_01624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05257__S1 (.I(_01624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05237__S1 (.I(_01624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05168__S1 (.I(_01624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05133__S1 (.I(_01624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05786__B (.I(_01626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05766__B (.I(_01626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05689__B (.I(_01626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05678__B (.I(_01626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05601__B (.I(_01626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05590__B (.I(_01626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05513__B (.I(_01626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05502__B (.I(_01626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05425__B (.I(_01626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05414__B (.I(_01626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05337__B (.I(_01626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05326__B (.I(_01626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05249__B (.I(_01626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05238__B (.I(_01626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05148__B (.I(_01626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05135__B (.I(_01626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05137__B2 (.I(_01627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05778__C (.I(_01628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05767__C (.I(_01628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05690__C (.I(_01628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05679__C (.I(_01628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05602__C (.I(_01628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05591__C (.I(_01628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05514__C (.I(_01628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05503__C (.I(_01628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05426__C (.I(_01628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05415__C (.I(_01628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05338__C (.I(_01628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05327__C (.I(_01628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05250__C (.I(_01628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05239__C (.I(_01628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05149__C (.I(_01628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05137__C (.I(_01628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05138__A3 (.I(_01629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05203__A2 (.I(_01631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05141__A2 (.I(_01632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05775__A1 (.I(_01636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05755__A1 (.I(_01636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05687__A1 (.I(_01636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05667__A1 (.I(_01636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05599__A1 (.I(_01636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05579__A1 (.I(_01636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05541__A1 (.I(_01636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05511__A1 (.I(_01636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05453__A1 (.I(_01636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05423__A1 (.I(_01636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05365__A1 (.I(_01636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05335__A1 (.I(_01636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05277__A1 (.I(_01636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05247__A1 (.I(_01636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05184__A1 (.I(_01636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05146__A1 (.I(_01636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05149__B1 (.I(_01638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05148__A2 (.I(_01639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05165__A2 (.I(_01641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05779__S1 (.I(_01642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05759__S1 (.I(_01642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05691__S1 (.I(_01642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05671__S1 (.I(_01642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05603__S1 (.I(_01642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05583__S1 (.I(_01642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05515__S1 (.I(_01642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05495__S1 (.I(_01642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05441__S1 (.I(_01642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05427__S1 (.I(_01642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05353__S1 (.I(_01642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05339__S1 (.I(_01642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05265__S1 (.I(_01642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05251__S1 (.I(_01642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05170__S1 (.I(_01642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05151__S1 (.I(_01642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05152__A2 (.I(_01643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05792__A1 (.I(_01645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05766__A1 (.I(_01645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05704__A1 (.I(_01645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05678__A1 (.I(_01645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05616__A1 (.I(_01645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05590__A1 (.I(_01645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05528__A1 (.I(_01645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05518__A1 (.I(_01645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05440__A1 (.I(_01645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05430__A1 (.I(_01645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05352__A1 (.I(_01645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05342__A1 (.I(_01645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05264__A1 (.I(_01645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05254__A1 (.I(_01645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05169__A1 (.I(_01645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05157__A1 (.I(_01645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05791__S0 (.I(_01646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05781__S0 (.I(_01646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05703__S0 (.I(_01646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05693__S0 (.I(_01646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05615__S0 (.I(_01646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05605__S0 (.I(_01646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05527__S0 (.I(_01646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05517__S0 (.I(_01646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05439__S0 (.I(_01646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05429__S0 (.I(_01646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05351__S0 (.I(_01646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05341__S0 (.I(_01646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05263__S0 (.I(_01646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05253__S0 (.I(_01646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05168__S0 (.I(_01646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05155__S0 (.I(_01646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05157__A2 (.I(_01647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05805__B (.I(_01648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05792__B (.I(_01648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05717__B (.I(_01648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05704__B (.I(_01648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05616__B (.I(_01648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05606__B (.I(_01648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05528__B (.I(_01648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05518__B (.I(_01648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05440__B (.I(_01648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05430__B (.I(_01648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05352__B (.I(_01648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05342__B (.I(_01648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05264__B (.I(_01648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05254__B (.I(_01648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05169__B (.I(_01648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05157__B (.I(_01648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05159__A2 (.I(_01650_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05800__S1 (.I(_01652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05795__S1 (.I(_01652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05712__S1 (.I(_01652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05707__S1 (.I(_01652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05624__S1 (.I(_01652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05619__S1 (.I(_01652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05536__S1 (.I(_01652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05531__S1 (.I(_01652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05448__S1 (.I(_01652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05443__S1 (.I(_01652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05360__S1 (.I(_01652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05355__S1 (.I(_01652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05272__S1 (.I(_01652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05267__S1 (.I(_01652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05172__S1 (.I(_01652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05161__S1 (.I(_01652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05801__B (.I(_01654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05796__B (.I(_01654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05708__B (.I(_01654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05698__B (.I(_01654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05620__B (.I(_01654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05610__B (.I(_01654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05532__B (.I(_01654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05522__B (.I(_01654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05444__B (.I(_01654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05434__B (.I(_01654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05356__B (.I(_01654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05346__B (.I(_01654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05268__B (.I(_01654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05258__B (.I(_01654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05173__B (.I(_01654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05163__B (.I(_01654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05164__B2 (.I(_01655_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05165__A3 (.I(_01656_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05187__A1 (.I(_01657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05169__A2 (.I(_01660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05173__A2 (.I(_01664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05186__A2 (.I(_01666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05799__A1 (.I(_01667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05715__A1 (.I(_01667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05711__A1 (.I(_01667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05627__A1 (.I(_01667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05623__A1 (.I(_01667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05539__A1 (.I(_01667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05535__A1 (.I(_01667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05451__A1 (.I(_01667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05447__A1 (.I(_01667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05363__A1 (.I(_01667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05359__A1 (.I(_01667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05275__A1 (.I(_01667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05271__A1 (.I(_01667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05192__I (.I(_01667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05182__A1 (.I(_01667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05178__A1 (.I(_01667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06135__A1 (.I(_01668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05798__S1 (.I(_01668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05734__S1 (.I(_01668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05710__S1 (.I(_01668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05622__S1 (.I(_01668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05534__S1 (.I(_01668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05450__S1 (.I(_01668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05446__S1 (.I(_01668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05362__S1 (.I(_01668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05358__S1 (.I(_01668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05274__S1 (.I(_01668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05270__S1 (.I(_01668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05196__I (.I(_01668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05189__I (.I(_01668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05181__S1 (.I(_01668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05177__S1 (.I(_01668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05178__A2 (.I(_01669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05185__A2 (.I(_01672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05182__A2 (.I(_01673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05186__A3 (.I(_01677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05202__A1 (.I(_01679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06493__A1 (.I(_01680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06492__A1 (.I(_01680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05811__S0 (.I(_01680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05723__S0 (.I(_01680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05635__S0 (.I(_01680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05633__S0 (.I(_01680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05547__S0 (.I(_01680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05545__S0 (.I(_01680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05459__S0 (.I(_01680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05457__S0 (.I(_01680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05371__S0 (.I(_01680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05369__S0 (.I(_01680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05283__S0 (.I(_01680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05281__S0 (.I(_01680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05193__S0 (.I(_01680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05190__S0 (.I(_01680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06496__A1 (.I(_01681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05811__S1 (.I(_01681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05723__S1 (.I(_01681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05721__S1 (.I(_01681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05635__S1 (.I(_01681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05633__S1 (.I(_01681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05547__S1 (.I(_01681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05545__S1 (.I(_01681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05459__S1 (.I(_01681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05457__S1 (.I(_01681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05371__S1 (.I(_01681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05369__S1 (.I(_01681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05283__S1 (.I(_01681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05281__S1 (.I(_01681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05193__S1 (.I(_01681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05190__S1 (.I(_01681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05191__A2 (.I(_01682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05816__A1 (.I(_01684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05812__A1 (.I(_01684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05728__A1 (.I(_01684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05724__A1 (.I(_01684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05640__A1 (.I(_01684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05636__A1 (.I(_01684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05552__A1 (.I(_01684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05548__A1 (.I(_01684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05464__A1 (.I(_01684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05460__A1 (.I(_01684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05376__A1 (.I(_01684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05372__A1 (.I(_01684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05288__A1 (.I(_01684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05284__A1 (.I(_01684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05200__A1 (.I(_01684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05194__A1 (.I(_01684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05815__S0 (.I(_01687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05809__S0 (.I(_01687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05727__S0 (.I(_01687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05721__S0 (.I(_01687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05639__S0 (.I(_01687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05637__S0 (.I(_01687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05551__S0 (.I(_01687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05549__S0 (.I(_01687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05463__S0 (.I(_01687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05461__S0 (.I(_01687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05375__S0 (.I(_01687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05373__S0 (.I(_01687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05287__S0 (.I(_01687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05285__S0 (.I(_01687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05199__S0 (.I(_01687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05197__S0 (.I(_01687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05815__S1 (.I(_01688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05809__S1 (.I(_01688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05727__S1 (.I(_01688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05725__S1 (.I(_01688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05639__S1 (.I(_01688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05637__S1 (.I(_01688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05551__S1 (.I(_01688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05549__S1 (.I(_01688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05463__S1 (.I(_01688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05461__S1 (.I(_01688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05375__S1 (.I(_01688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05373__S1 (.I(_01688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05287__S1 (.I(_01688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05285__S1 (.I(_01688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05199__S1 (.I(_01688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05197__S1 (.I(_01688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05200__A2 (.I(_01691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05202__A2 (.I(_01693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05205__A2 (.I(_01695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05207__A2 (.I(_01697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05209__A2 (.I(_01699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05241__A2 (.I(_01703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05214__A2 (.I(_01704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05216__A2 (.I(_01706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05218__A2 (.I(_01708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05220__A2 (.I(_01710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05223__A2 (.I(_01713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05225__A2 (.I(_01715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05227__A2 (.I(_01717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05229__A2 (.I(_01719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05232__A2 (.I(_01722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05234__A2 (.I(_01724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05239__A2 (.I(_01725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05238__A2 (.I(_01728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05239__B2 (.I(_01729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05240__A3 (.I(_01730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05291__A2 (.I(_01732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05243__A2 (.I(_01733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05247__A2 (.I(_01737_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05250__B1 (.I(_01738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05249__A2 (.I(_01739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05260__A2 (.I(_01741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05252__A2 (.I(_01742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05254__A2 (.I(_01744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05256__A2 (.I(_01746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05260__A3 (.I(_01750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05280__A1 (.I(_01751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05264__A2 (.I(_01754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05268__A2 (.I(_01758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05279__A2 (.I(_01760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05271__A2 (.I(_01761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05278__A2 (.I(_01764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05275__A2 (.I(_01765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05279__A3 (.I(_01769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05290__A1 (.I(_01771_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05282__A2 (.I(_01772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05288__A2 (.I(_01778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05290__A2 (.I(_01780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05293__A2 (.I(_01782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05295__A2 (.I(_01784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05297__A2 (.I(_01786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05329__A2 (.I(_01790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05309__A1 (.I(_01792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05304__A2 (.I(_01793_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05308__A2 (.I(_01797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05329__A3 (.I(_01799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05311__A2 (.I(_01800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05313__A2 (.I(_01802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05315__A2 (.I(_01804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05317__A2 (.I(_01806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05320__A2 (.I(_01809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05322__A2 (.I(_01811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05324__A2 (.I(_01813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05326__A2 (.I(_01815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05327__B2 (.I(_01816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05328__A3 (.I(_01817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05379__A2 (.I(_01819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05331__A2 (.I(_01820_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05338__B1 (.I(_01825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05348__A2 (.I(_01828_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05340__A2 (.I(_01829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05346__A2 (.I(_01835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05347__B2 (.I(_01836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05348__A3 (.I(_01837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05368__A1 (.I(_01838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05357__A2 (.I(_01842_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05356__A2 (.I(_01845_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05367__A2 (.I(_01847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05359__A2 (.I(_01848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05366__A2 (.I(_01851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05363__A2 (.I(_01852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05367__A3 (.I(_01856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05378__A1 (.I(_01858_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05370__A2 (.I(_01859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05376__A2 (.I(_01865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05378__A2 (.I(_01867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05381__A2 (.I(_01869_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05383__A2 (.I(_01871_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05385__A2 (.I(_01873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05417__A2 (.I(_01877_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05390__A2 (.I(_01878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05392__A2 (.I(_01880_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05397__A2 (.I(_01881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05396__A2 (.I(_01884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05417__A3 (.I(_01886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05401__A2 (.I(_01889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05403__A2 (.I(_01891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05405__A2 (.I(_01893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05408__A2 (.I(_01896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05410__A2 (.I(_01898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05414__A2 (.I(_01902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05416__A3 (.I(_01904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05467__A2 (.I(_01906_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05419__A2 (.I(_01907_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05423__A2 (.I(_01911_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05426__B1 (.I(_01912_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05436__A2 (.I(_01915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05428__A2 (.I(_01916_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05430__A2 (.I(_01918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05432__A2 (.I(_01920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05436__A3 (.I(_01924_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05456__A1 (.I(_01925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05440__A2 (.I(_01928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05445__A2 (.I(_01929_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05444__A2 (.I(_01932_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05455__A2 (.I(_01934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05447__A2 (.I(_01935_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05454__A2 (.I(_01938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05451__A2 (.I(_01939_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05455__A3 (.I(_01943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05466__A1 (.I(_01945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05458__A2 (.I(_01946_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05464__A2 (.I(_01952_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05466__A2 (.I(_01954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05469__A2 (.I(_01956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05471__A2 (.I(_01958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05473__A2 (.I(_01960_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05505__A2 (.I(_01964_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05484__A2 (.I(_01971_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05505__A3 (.I(_01973_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05489__A2 (.I(_01976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05491__A2 (.I(_01978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05493__A2 (.I(_01980_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05496__A2 (.I(_01983_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05498__A2 (.I(_01985_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05502__A2 (.I(_01989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05504__A3 (.I(_01991_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05555__A2 (.I(_01993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05507__A2 (.I(_01994_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05514__B1 (.I(_01999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05513__A2 (.I(_02000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05524__A2 (.I(_02002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05516__A2 (.I(_02003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05518__A2 (.I(_02005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05520__A2 (.I(_02007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05523__B2 (.I(_02010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05524__A3 (.I(_02011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05544__A1 (.I(_02012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05526__A2 (.I(_02013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05528__A2 (.I(_02015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05532__A2 (.I(_02019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05543__A2 (.I(_02021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05535__A2 (.I(_02022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05542__A2 (.I(_02025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05539__A2 (.I(_02026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05543__A3 (.I(_02030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05554__A1 (.I(_02032_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05546__A2 (.I(_02033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05552__A2 (.I(_02039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05554__A2 (.I(_02041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05557__A2 (.I(_02043_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05561__A2 (.I(_02047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05593__A2 (.I(_02051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05568__A2 (.I(_02054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05573__A2 (.I(_02055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05572__A2 (.I(_02058_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05593__A3 (.I(_02060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05575__A2 (.I(_02061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05577__A2 (.I(_02063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05582__A2 (.I(_02064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05579__A2 (.I(_02065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05581__A2 (.I(_02067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05584__A2 (.I(_02070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05586__A2 (.I(_02072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05591__A2 (.I(_02073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05590__A2 (.I(_02076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05591__B2 (.I(_02077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05592__A3 (.I(_02078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05643__A2 (.I(_02080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05595__A2 (.I(_02081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05597__A2 (.I(_02083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05599__A2 (.I(_02085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05602__B1 (.I(_02086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05601__A2 (.I(_02087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05612__A2 (.I(_02089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05604__A2 (.I(_02090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05611__A1 (.I(_02091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05606__A2 (.I(_02092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05608__A2 (.I(_02094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05611__B1 (.I(_02095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05612__A3 (.I(_02098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05632__A1 (.I(_02099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05616__A2 (.I(_02102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05618__A2 (.I(_02104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05620__A2 (.I(_02106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05631__A2 (.I(_02108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05623__A2 (.I(_02109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05630__A2 (.I(_02112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05627__A2 (.I(_02113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05631__A3 (.I(_02117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05642__A1 (.I(_02119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05634__A2 (.I(_02120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05636__A2 (.I(_02122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05640__A2 (.I(_02126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05642__A2 (.I(_02128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05643__B (.I(_02129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05645__A2 (.I(_02130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05649__A2 (.I(_02134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05681__A2 (.I(_02138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05661__A2 (.I(_02142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05658__A2 (.I(_02143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05660__A2 (.I(_02145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05681__A3 (.I(_02147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05663__A2 (.I(_02148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05665__A2 (.I(_02150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05670__A2 (.I(_02151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05667__A2 (.I(_02152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05669__A2 (.I(_02154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05672__A2 (.I(_02157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05680__A3 (.I(_02165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05731__A2 (.I(_02167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05683__A2 (.I(_02168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05685__A2 (.I(_02170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05690__B1 (.I(_02173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05700__A2 (.I(_02176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05692__A2 (.I(_02177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05699__A1 (.I(_02178_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05696__A2 (.I(_02181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05700__A3 (.I(_02185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05720__A1 (.I(_02186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05709__A2 (.I(_02190_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05706__A2 (.I(_02191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05708__A2 (.I(_02193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05719__A2 (.I(_02195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05711__A2 (.I(_02196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05718__A2 (.I(_02199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05715__A2 (.I(_02200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05719__A3 (.I(_02204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05730__A1 (.I(_02206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05722__A2 (.I(_02207_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05724__A2 (.I(_02209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05728__A2 (.I(_02213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05730__A2 (.I(_02215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05733__A2 (.I(_02217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05740__A2 (.I(_02220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05737__A2 (.I(_02221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05769__A2 (.I(_02225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05746__A2 (.I(_02230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05748__A2 (.I(_02232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05769__A3 (.I(_02234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05753__A2 (.I(_02237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05755__A2 (.I(_02239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05757__A2 (.I(_02241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05758__B2 (.I(_02242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05760__A2 (.I(_02244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05762__A2 (.I(_02246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05767__B2 (.I(_02251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05768__A3 (.I(_02252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05771__A2 (.I(_02255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05775__A2 (.I(_02259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05777__A2 (.I(_02261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05788__A2 (.I(_02263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05780__A2 (.I(_02264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05782__A2 (.I(_02266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05787__B2 (.I(_02271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05788__A3 (.I(_02272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05808__A1 (.I(_02273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05797__A2 (.I(_02277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05797__B1 (.I(_02279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05796__A2 (.I(_02280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05807__A2 (.I(_02282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05799__A2 (.I(_02283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05803__A2 (.I(_02287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05806__B1 (.I(_02288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05807__A3 (.I(_02291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05818__A1 (.I(_02293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05810__A2 (.I(_02294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05817__B1 (.I(_02299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05816__A2 (.I(_02300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05818__A2 (.I(_02302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09361__A1 (.I(_02305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08654__A1 (.I(_02305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08458__A2 (.I(_02305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08447__A1 (.I(_02305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08443__A2 (.I(_02305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08404__A1 (.I(_02305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08373__A1 (.I(_02305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08334__B (.I(_02305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08007__A1 (.I(_02305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05985__A1 (.I(_02305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05884__A1 (.I(_02305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05862__A1 (.I(_02305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05846__A1 (.I(_02305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05845__A1 (.I(_02305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09369__A2 (.I(_02306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08226__A1 (.I(_02306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05992__A1 (.I(_02306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05970__I (.I(_02306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05920__A2 (.I(_02306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05841__S (.I(_02306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05832__A1 (.I(_02306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05831__A1 (.I(_02306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05824__A1 (.I(_02306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07733__A1 (.I(_02309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05977__A1 (.I(_02309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05974__A1 (.I(_02309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05876__A1 (.I(_02309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05870__A1 (.I(_02309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05869__A1 (.I(_02309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05848__A2 (.I(_02309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05843__A1 (.I(_02309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05826__A1 (.I(_02309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09380__A1 (.I(_02311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09360__A1 (.I(_02311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08523__A1 (.I(_02311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07682__A2 (.I(_02311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07671__A1 (.I(_02311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06474__A1 (.I(_02311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05913__A1 (.I(_02311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05912__A1 (.I(_02311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05859__A1 (.I(_02311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05835__A1 (.I(_02311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05834__A1 (.I(_02311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08803__A1 (.I(_02312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06001__A1 (.I(_02312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05831__A2 (.I(_02312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08424__A2 (.I(_02313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08372__A2 (.I(_02313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08334__A2 (.I(_02313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07741__A1 (.I(_02313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05992__A2 (.I(_02313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05975__A2 (.I(_02313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05919__A2 (.I(_02313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05910__A2 (.I(_02313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05901__I (.I(_02313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05900__A2 (.I(_02313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05881__A2 (.I(_02313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05830__A3 (.I(_02313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09563__A2 (.I(_02320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05949__A1 (.I(_02320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05948__A1 (.I(_02320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05946__A1 (.I(_02320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05945__A1 (.I(_02320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05943__A1 (.I(_02320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05942__A1 (.I(_02320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05940__A1 (.I(_02320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05939__A1 (.I(_02320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05937__A1 (.I(_02320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05936__A1 (.I(_02320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05934__A1 (.I(_02320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05933__A1 (.I(_02320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05840__A1 (.I(_02320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05839__A2 (.I(_02320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09565__A1 (.I(_02321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09563__A1 (.I(_02321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05947__A1 (.I(_02321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05944__A1 (.I(_02321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05941__A1 (.I(_02321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05938__A1 (.I(_02321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05935__A1 (.I(_02321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05932__A1 (.I(_02321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05838__A2 (.I(_02321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08725__A1 (.I(_02324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05864__A2 (.I(_02324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05841__I1 (.I(_02324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08120__B2 (.I(_02325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07734__A1 (.I(_02325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05877__A3 (.I(_02325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05870__A2 (.I(_02325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05869__A2 (.I(_02325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05842__A2 (.I(_02325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08247__A1 (.I(_02332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07737__A2 (.I(_02332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06476__A2 (.I(_02332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05998__B (.I(_02332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05997__B (.I(_02332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05996__B (.I(_02332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05965__A1 (.I(_02332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05903__A1 (.I(_02332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05851__A1 (.I(_02332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08240__A1 (.I(_02333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07740__A1 (.I(_02333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05852__B (.I(_02333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05851__A2 (.I(_02333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09386__A4 (.I(_02337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08288__A1 (.I(_02337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05857__A1 (.I(_02337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09361__A3 (.I(_02338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08628__B (.I(_02338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05897__A1 (.I(_02338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05874__A2 (.I(_02338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05863__A2 (.I(_02338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05859__B (.I(_02338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05857__A3 (.I(_02338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09387__A1 (.I(_02339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05857__A4 (.I(_02339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09368__A1 (.I(_02341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05863__A1 (.I(_02341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08722__A1 (.I(_02343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08276__A1 (.I(_02343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05861__A1 (.I(_02343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09380__A2 (.I(_02344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09361__A2 (.I(_02344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05862__A2 (.I(_02344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09390__A2 (.I(_02348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09388__A1 (.I(_02348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05866__A2 (.I(_02348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08725__A2 (.I(_02356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07738__A2 (.I(_02356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05976__A2 (.I(_02356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05925__A2 (.I(_02356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05875__A3 (.I(_02356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08631__A1 (.I(_02361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05965__B2 (.I(_02361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05918__A1 (.I(_02361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05891__A1 (.I(_02361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08629__A1 (.I(_02372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08619__S (.I(_02372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08586__I (.I(_02372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05980__I (.I(_02372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05918__A3 (.I(_02372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05891__A2 (.I(_02372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08724__I0 (.I(_02381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05909__A1 (.I(_02381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08446__A2 (.I(_02391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05926__A2 (.I(_02391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05915__A2 (.I(_02391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08625__A2 (.I(_02394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05979__A2 (.I(_02394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05917__A1 (.I(_02394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07743__A2 (.I(_02395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05916__A2 (.I(_02395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05982__A3 (.I(_02401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05921__A2 (.I(_02401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08724__I1 (.I(_02406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05928__A2 (.I(_02406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05926__A3 (.I(_02406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05931__I (.I(_02411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08635__A1 (.I(_02431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05998__A1 (.I(_02431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05997__A2 (.I(_02431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05965__A2 (.I(_02431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08800__A1 (.I(_02433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08563__A1 (.I(_02433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08562__A2 (.I(_02433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08442__A1 (.I(_02433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07685__B (.I(_02433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06487__A3 (.I(_02433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05994__B (.I(_02433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05990__A2 (.I(_02433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05968__A2 (.I(_02433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08372__A1 (.I(_02436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08334__A1 (.I(_02436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05971__A1 (.I(_02436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08427__A2 (.I(_02438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08426__C (.I(_02438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05977__A3 (.I(_02438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05974__A4 (.I(_02438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08627__B2 (.I(_02445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08624__B (.I(_02445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08623__A2 (.I(_02445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08622__A2 (.I(_02445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08584__S (.I(_02445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08582__S (.I(_02445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08580__S (.I(_02445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08578__S (.I(_02445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08576__S (.I(_02445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08574__S (.I(_02445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08572__S (.I(_02445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08570__S (.I(_02445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08568__S (.I(_02445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08566__S (.I(_02445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08564__S (.I(_02445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05981__B (.I(_02445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08654__A2 (.I(_02448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08632__A2 (.I(_02448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08624__A2 (.I(_02448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08523__A2 (.I(_02448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06474__A2 (.I(_02448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05993__C (.I(_02448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05985__A2 (.I(_02448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08800__A2 (.I(_02453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05993__B (.I(_02453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06188__S (.I(_02460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06065__A1 (.I(_02460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06059__A1 (.I(_02460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06053__A1 (.I(_02460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06047__A1 (.I(_02460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06041__A1 (.I(_02460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06035__A1 (.I(_02460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06029__A1 (.I(_02460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06023__A2 (.I(_02460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06005__A1 (.I(_02460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06004__A2 (.I(_02460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09488__A1 (.I(_02469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08765__A1 (.I(_02469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08289__A1 (.I(_02469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07783__A1 (.I(_02469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07448__A1 (.I(_02469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06735__A1 (.I(_02469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06426__A1 (.I(_02469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06117__A1 (.I(_02469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06019__A1 (.I(_02469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06018__I (.I(_02474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09524__A1 (.I(_02475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09342__A1 (.I(_02475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09324__A1 (.I(_02475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09288__A1 (.I(_02475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09252__A1 (.I(_02475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09192__A1 (.I(_02475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09137__A1 (.I(_02475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08883__A1 (.I(_02475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08858__A1 (.I(_02475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08782__A1 (.I(_02475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07747__A1 (.I(_02475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07710__A1 (.I(_02475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07692__A1 (.I(_02475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06212__A1 (.I(_02475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06099__A1 (.I(_02475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06019__A2 (.I(_02475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06069__A1 (.I(_02477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06068__A2 (.I(_02477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06063__A1 (.I(_02477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06062__A2 (.I(_02477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06057__A1 (.I(_02477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06056__A2 (.I(_02477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06051__A1 (.I(_02477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06050__A2 (.I(_02477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06045__A1 (.I(_02477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06044__A2 (.I(_02477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06039__A1 (.I(_02477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06038__A2 (.I(_02477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06033__A1 (.I(_02477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06032__A2 (.I(_02477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06027__A1 (.I(_02477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06026__A2 (.I(_02477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06184__S (.I(_02478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06180__S (.I(_02478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06176__S (.I(_02478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06172__S (.I(_02478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06168__S (.I(_02478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06164__S (.I(_02478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06159__A1 (.I(_02478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06155__S (.I(_02478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06064__A1 (.I(_02478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06058__A1 (.I(_02478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06052__A1 (.I(_02478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06046__A1 (.I(_02478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06040__A1 (.I(_02478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06034__A1 (.I(_02478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06028__A1 (.I(_02478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06022__A2 (.I(_02478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09191__I (.I(_02481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08857__I (.I(_02481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07819__I (.I(_02481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07483__I (.I(_02481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07153__I (.I(_02481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06789__I (.I(_02481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06425__I (.I(_02481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06025__I (.I(_02481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06410__A1 (.I(_02482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06391__A1 (.I(_02482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06373__A1 (.I(_02482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06354__A1 (.I(_02482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06335__A1 (.I(_02482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06314__A1 (.I(_02482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06295__A1 (.I(_02482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06276__A1 (.I(_02482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06258__A1 (.I(_02482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06237__A1 (.I(_02482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06215__A1 (.I(_02482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06140__A1 (.I(_02482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06120__A1 (.I(_02482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06102__A1 (.I(_02482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06083__A1 (.I(_02482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06027__A2 (.I(_02482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09196__I (.I(_02486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08862__I (.I(_02486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07824__I (.I(_02486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07488__I (.I(_02486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07158__I (.I(_02486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06794__I (.I(_02486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06430__I (.I(_02486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06031__I (.I(_02486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06412__A1 (.I(_02487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06393__A1 (.I(_02487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06375__A1 (.I(_02487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06356__A1 (.I(_02487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06337__A1 (.I(_02487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06316__A1 (.I(_02487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06297__A1 (.I(_02487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06278__A1 (.I(_02487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06260__A1 (.I(_02487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06239__A1 (.I(_02487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06217__A1 (.I(_02487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06142__A1 (.I(_02487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06122__A1 (.I(_02487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06104__A1 (.I(_02487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06085__A1 (.I(_02487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06033__A2 (.I(_02487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09199__I (.I(_02491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08865__I (.I(_02491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07827__I (.I(_02491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07491__I (.I(_02491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07161__I (.I(_02491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06797__I (.I(_02491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06433__I (.I(_02491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06037__I (.I(_02491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06414__A1 (.I(_02492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06395__A1 (.I(_02492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06377__A1 (.I(_02492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06358__A1 (.I(_02492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06339__A1 (.I(_02492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06318__A1 (.I(_02492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06299__A1 (.I(_02492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06280__A1 (.I(_02492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06262__A1 (.I(_02492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06241__A1 (.I(_02492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06219__A1 (.I(_02492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06144__A1 (.I(_02492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06124__A1 (.I(_02492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06106__A1 (.I(_02492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06087__A1 (.I(_02492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06039__A2 (.I(_02492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09202__I (.I(_02496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08868__I (.I(_02496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07830__I (.I(_02496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07494__I (.I(_02496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07164__I (.I(_02496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06800__I (.I(_02496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06436__I (.I(_02496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06043__I (.I(_02496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06416__A1 (.I(_02497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06397__A1 (.I(_02497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06379__A1 (.I(_02497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06360__A1 (.I(_02497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06341__A1 (.I(_02497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06320__A1 (.I(_02497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06301__A1 (.I(_02497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06282__A1 (.I(_02497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06264__A1 (.I(_02497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06243__A1 (.I(_02497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06221__A1 (.I(_02497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06146__A1 (.I(_02497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06126__A1 (.I(_02497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06108__A1 (.I(_02497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06089__A1 (.I(_02497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06045__A2 (.I(_02497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09205__I (.I(_02501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08871__I (.I(_02501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07833__I (.I(_02501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07497__I (.I(_02501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07167__I (.I(_02501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06803__I (.I(_02501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06439__I (.I(_02501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06049__I (.I(_02501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06418__A1 (.I(_02502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06399__A1 (.I(_02502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06381__A1 (.I(_02502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06362__A1 (.I(_02502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06343__A1 (.I(_02502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06322__A1 (.I(_02502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06303__A1 (.I(_02502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06284__A1 (.I(_02502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06266__A1 (.I(_02502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06245__A1 (.I(_02502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06223__A1 (.I(_02502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06148__A1 (.I(_02502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06128__A1 (.I(_02502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06110__A1 (.I(_02502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06091__A1 (.I(_02502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06051__A2 (.I(_02502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09208__I (.I(_02506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08874__I (.I(_02506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07836__I (.I(_02506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07500__I (.I(_02506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07170__I (.I(_02506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06806__I (.I(_02506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06442__I (.I(_02506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06055__I (.I(_02506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06420__A1 (.I(_02507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06401__A1 (.I(_02507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06383__A1 (.I(_02507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06364__A1 (.I(_02507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06345__A1 (.I(_02507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06324__A1 (.I(_02507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06305__A1 (.I(_02507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06286__A1 (.I(_02507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06268__A1 (.I(_02507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06247__A1 (.I(_02507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06225__A1 (.I(_02507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06150__A1 (.I(_02507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06130__A1 (.I(_02507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06112__A1 (.I(_02507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06093__A1 (.I(_02507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06057__A2 (.I(_02507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09211__I (.I(_02511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08877__I (.I(_02511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07839__I (.I(_02511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07503__I (.I(_02511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07173__I (.I(_02511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06809__I (.I(_02511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06445__I (.I(_02511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06061__I (.I(_02511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06422__A1 (.I(_02512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06403__A1 (.I(_02512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06385__A1 (.I(_02512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06366__A1 (.I(_02512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06347__A1 (.I(_02512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06326__A1 (.I(_02512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06307__A1 (.I(_02512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06288__A1 (.I(_02512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06270__A1 (.I(_02512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06249__A1 (.I(_02512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06227__A1 (.I(_02512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06152__A1 (.I(_02512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06132__A1 (.I(_02512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06114__A1 (.I(_02512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06095__A1 (.I(_02512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06063__A2 (.I(_02512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09214__I (.I(_02516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08880__I (.I(_02516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07842__I (.I(_02516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07506__I (.I(_02516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07176__I (.I(_02516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06812__I (.I(_02516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06448__I (.I(_02516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06067__I (.I(_02516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06424__A1 (.I(_02517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06405__A1 (.I(_02517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06387__A1 (.I(_02517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06368__A1 (.I(_02517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06349__A1 (.I(_02517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06328__A1 (.I(_02517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06309__A1 (.I(_02517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06290__A1 (.I(_02517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06272__A1 (.I(_02517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06251__A1 (.I(_02517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06229__A1 (.I(_02517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06154__A1 (.I(_02517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06134__A1 (.I(_02517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06116__A1 (.I(_02517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06097__A1 (.I(_02517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06069__A2 (.I(_02517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09252__A2 (.I(_02524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09173__A1 (.I(_02524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08975__A1 (.I(_02524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07801__A1 (.I(_02524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07635__A1 (.I(_02524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07394__A1 (.I(_02524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07012__A1 (.I(_02524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06905__A1 (.I(_02524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06080__A1 (.I(_02524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06079__I (.I(_02527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09542__A1 (.I(_02528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09453__A1 (.I(_02528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09435__A1 (.I(_02528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09417__A1 (.I(_02528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09399__A1 (.I(_02528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08924__A1 (.I(_02528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08636__A1 (.I(_02528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08544__A1 (.I(_02528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07484__A1 (.I(_02528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06887__A1 (.I(_02528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06790__A1 (.I(_02528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06516__A1 (.I(_02528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06498__A1 (.I(_02528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06137__A1 (.I(_02528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06117__A2 (.I(_02528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06080__A2 (.I(_02528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06097__A2 (.I(_02530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06096__A2 (.I(_02530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06095__A2 (.I(_02530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06094__A2 (.I(_02530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06093__A2 (.I(_02530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06092__A2 (.I(_02530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06091__A2 (.I(_02530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06090__A2 (.I(_02530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06089__A2 (.I(_02530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06088__A2 (.I(_02530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06087__A2 (.I(_02530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06086__A2 (.I(_02530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06085__A2 (.I(_02530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06084__A2 (.I(_02530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06083__A2 (.I(_02530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06082__A2 (.I(_02530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08839__A1 (.I(_02539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08122__A1 (.I(_02539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07987__A1 (.I(_02539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07322__A1 (.I(_02539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06753__A1 (.I(_02539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06573__A1 (.I(_02539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06516__A2 (.I(_02539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06161__A1 (.I(_02539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06099__A2 (.I(_02539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06116__A2 (.I(_02541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06115__A2 (.I(_02541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06114__A2 (.I(_02541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06113__A2 (.I(_02541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06112__A2 (.I(_02541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06111__A2 (.I(_02541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06110__A2 (.I(_02541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06109__A2 (.I(_02541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06108__A2 (.I(_02541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06107__A2 (.I(_02541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06106__A2 (.I(_02541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06105__A2 (.I(_02541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06104__A2 (.I(_02541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06103__A2 (.I(_02541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06102__A2 (.I(_02541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06101__A2 (.I(_02541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06134__A2 (.I(_02551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06133__A2 (.I(_02551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06132__A2 (.I(_02551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06131__A2 (.I(_02551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06130__A2 (.I(_02551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06129__A2 (.I(_02551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06128__A2 (.I(_02551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06127__A2 (.I(_02551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06126__A2 (.I(_02551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06125__A2 (.I(_02551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06124__A2 (.I(_02551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06123__A2 (.I(_02551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06122__A2 (.I(_02551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06121__A2 (.I(_02551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06120__A2 (.I(_02551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06119__A2 (.I(_02551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09506__A1 (.I(_02561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09192__A2 (.I(_02561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07969__A1 (.I(_02561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07653__A1 (.I(_02561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07412__A1 (.I(_02561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07030__A1 (.I(_02561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06699__A1 (.I(_02561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06451__A1 (.I(_02561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06137__A2 (.I(_02561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06154__A2 (.I(_02563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06153__A2 (.I(_02563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06152__A2 (.I(_02563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06151__A2 (.I(_02563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06150__A2 (.I(_02563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06149__A2 (.I(_02563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06148__A2 (.I(_02563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06147__A2 (.I(_02563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06146__A2 (.I(_02563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06145__A2 (.I(_02563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06144__A2 (.I(_02563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06143__A2 (.I(_02563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06142__A2 (.I(_02563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06141__A2 (.I(_02563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06140__A2 (.I(_02563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06139__A2 (.I(_02563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09472__I0 (.I(_02573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09236__I0 (.I(_02573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08766__I0 (.I(_02573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08749__I0 (.I(_02573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07899__I0 (.I(_02573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07882__I0 (.I(_02573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07467__I0 (.I(_02573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07252__I0 (.I(_02573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07137__I0 (.I(_02573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07066__I0 (.I(_02573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07049__I0 (.I(_02573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06906__I0 (.I(_02573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06683__I0 (.I(_02573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06452__I0 (.I(_02573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06195__I0 (.I(_02573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06162__I0 (.I(_02573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06160__I (.I(_02576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09471__A1 (.I(_02577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09235__A1 (.I(_02577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08765__A2 (.I(_02577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08748__A1 (.I(_02577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07898__A1 (.I(_02577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07881__A1 (.I(_02577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07466__A1 (.I(_02577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07251__A1 (.I(_02577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07136__A1 (.I(_02577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07065__A1 (.I(_02577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07048__A1 (.I(_02577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06905__A2 (.I(_02577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06682__A1 (.I(_02577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06451__A2 (.I(_02577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06194__A1 (.I(_02577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06161__A2 (.I(_02577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06190__S (.I(_02578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06186__S (.I(_02578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06182__S (.I(_02578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06178__S (.I(_02578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06174__S (.I(_02578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06170__S (.I(_02578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06166__S (.I(_02578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06162__S (.I(_02578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09474__I0 (.I(_02581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09238__I0 (.I(_02581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08768__I0 (.I(_02581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08751__I0 (.I(_02581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07901__I0 (.I(_02581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07884__I0 (.I(_02581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07469__I0 (.I(_02581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07254__I0 (.I(_02581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07139__I0 (.I(_02581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07068__I0 (.I(_02581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07051__I0 (.I(_02581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06908__I0 (.I(_02581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06685__I0 (.I(_02581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06454__I0 (.I(_02581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06197__I0 (.I(_02581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06166__I0 (.I(_02581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09476__I0 (.I(_02584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09240__I0 (.I(_02584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08770__I0 (.I(_02584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08753__I0 (.I(_02584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07903__I0 (.I(_02584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07886__I0 (.I(_02584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07471__I0 (.I(_02584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07256__I0 (.I(_02584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07141__I0 (.I(_02584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07070__I0 (.I(_02584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07053__I0 (.I(_02584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06910__I0 (.I(_02584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06687__I0 (.I(_02584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06456__I0 (.I(_02584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06199__I0 (.I(_02584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06170__I0 (.I(_02584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09478__I0 (.I(_02587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09242__I0 (.I(_02587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08772__I0 (.I(_02587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08755__I0 (.I(_02587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07905__I0 (.I(_02587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07888__I0 (.I(_02587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07473__I0 (.I(_02587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07258__I0 (.I(_02587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07143__I0 (.I(_02587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07072__I0 (.I(_02587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07055__I0 (.I(_02587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06912__I0 (.I(_02587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06689__I0 (.I(_02587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06458__I0 (.I(_02587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06201__I0 (.I(_02587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06174__I0 (.I(_02587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09480__I0 (.I(_02590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09244__I0 (.I(_02590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08774__I0 (.I(_02590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08757__I0 (.I(_02590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07907__I0 (.I(_02590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07890__I0 (.I(_02590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07475__I0 (.I(_02590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07260__I0 (.I(_02590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07145__I0 (.I(_02590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07074__I0 (.I(_02590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07057__I0 (.I(_02590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06914__I0 (.I(_02590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06691__I0 (.I(_02590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06460__I0 (.I(_02590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06203__I0 (.I(_02590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06178__I0 (.I(_02590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09482__I0 (.I(_02593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09246__I0 (.I(_02593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08776__I0 (.I(_02593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08759__I0 (.I(_02593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07909__I0 (.I(_02593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07892__I0 (.I(_02593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07477__I0 (.I(_02593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07262__I0 (.I(_02593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07147__I0 (.I(_02593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07076__I0 (.I(_02593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07059__I0 (.I(_02593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06916__I0 (.I(_02593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06693__I0 (.I(_02593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06462__I0 (.I(_02593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06205__I0 (.I(_02593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06182__I0 (.I(_02593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09484__I0 (.I(_02596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09248__I0 (.I(_02596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08778__I0 (.I(_02596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08761__I0 (.I(_02596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07911__I0 (.I(_02596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07894__I0 (.I(_02596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07479__I0 (.I(_02596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07264__I0 (.I(_02596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07149__I0 (.I(_02596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07078__I0 (.I(_02596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07061__I0 (.I(_02596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06918__I0 (.I(_02596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06695__I0 (.I(_02596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06464__I0 (.I(_02596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06207__I0 (.I(_02596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06186__I0 (.I(_02596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09486__I0 (.I(_02599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09250__I0 (.I(_02599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08780__I0 (.I(_02599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08763__I0 (.I(_02599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07913__I0 (.I(_02599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07896__I0 (.I(_02599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07481__I0 (.I(_02599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07266__I0 (.I(_02599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07151__I0 (.I(_02599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07080__I0 (.I(_02599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07063__I0 (.I(_02599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06920__I0 (.I(_02599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06697__I0 (.I(_02599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06466__I0 (.I(_02599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06209__I0 (.I(_02599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06190__I0 (.I(_02599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09542__A2 (.I(_02602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09324__A2 (.I(_02602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09011__A1 (.I(_02602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07358__A1 (.I(_02602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07286__A1 (.I(_02602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07197__A1 (.I(_02602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06976__A1 (.I(_02602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06554__A1 (.I(_02602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06194__A2 (.I(_02602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06209__S (.I(_02603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06207__S (.I(_02603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06205__S (.I(_02603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06203__S (.I(_02603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06201__S (.I(_02603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06199__S (.I(_02603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06197__S (.I(_02603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06195__S (.I(_02603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09471__A2 (.I(_02612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08901__A1 (.I(_02612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08526__A1 (.I(_02612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07915__A1 (.I(_02612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07509__A1 (.I(_02612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06771__A1 (.I(_02612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06498__A2 (.I(_02612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06388__A1 (.I(_02612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06212__A2 (.I(_02612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06229__A2 (.I(_02614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06228__A2 (.I(_02614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06227__A2 (.I(_02614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06226__A2 (.I(_02614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06225__A2 (.I(_02614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06224__A2 (.I(_02614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06223__A2 (.I(_02614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06222__A2 (.I(_02614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06221__A2 (.I(_02614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06220__A2 (.I(_02614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06219__A2 (.I(_02614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06218__A2 (.I(_02614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06217__A2 (.I(_02614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06216__A2 (.I(_02614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06215__A2 (.I(_02614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06214__A2 (.I(_02614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09270__A1 (.I(_02625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08858__A2 (.I(_02625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08636__A2 (.I(_02625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07545__A1 (.I(_02625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07251__A2 (.I(_02625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07082__A1 (.I(_02625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06833__A1 (.I(_02625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06273__A1 (.I(_02625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06234__A1 (.I(_02625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09173__A2 (.I(_02626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09065__A1 (.I(_02626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07215__A1 (.I(_02626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07197__A2 (.I(_02626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07179__A1 (.I(_02626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07154__A1 (.I(_02626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06771__A2 (.I(_02626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06753__A2 (.I(_02626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06735__A2 (.I(_02626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06717__A1 (.I(_02626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06699__A2 (.I(_02626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06663__A1 (.I(_02626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06645__A1 (.I(_02626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06627__A1 (.I(_02626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06609__A1 (.I(_02626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06234__A2 (.I(_02626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06251__A2 (.I(_02628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06250__A2 (.I(_02628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06249__A2 (.I(_02628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06248__A2 (.I(_02628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06247__A2 (.I(_02628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06246__A2 (.I(_02628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06245__A2 (.I(_02628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06244__A2 (.I(_02628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06243__A2 (.I(_02628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06242__A2 (.I(_02628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06241__A2 (.I(_02628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06240__A2 (.I(_02628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06239__A2 (.I(_02628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06238__A2 (.I(_02628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06237__A2 (.I(_02628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06236__A2 (.I(_02628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09417__A2 (.I(_02638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09235__A2 (.I(_02638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09101__A1 (.I(_02638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07933__A1 (.I(_02638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07710__A2 (.I(_02638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07268__A1 (.I(_02638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06922__A1 (.I(_02638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06627__A2 (.I(_02638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06255__A1 (.I(_02638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08526__A2 (.I(_02639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07987__A2 (.I(_02639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07783__A2 (.I(_02639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07765__A1 (.I(_02639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07653__A2 (.I(_02639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07635__A2 (.I(_02639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07617__A1 (.I(_02639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07286__A2 (.I(_02639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06535__A1 (.I(_02639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06407__A1 (.I(_02639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06370__A1 (.I(_02639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06351__A1 (.I(_02639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06311__A1 (.I(_02639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06292__A1 (.I(_02639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06273__A2 (.I(_02639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06255__A2 (.I(_02639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06272__A2 (.I(_02641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06271__A2 (.I(_02641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06270__A2 (.I(_02641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06269__A2 (.I(_02641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06268__A2 (.I(_02641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06267__A2 (.I(_02641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06266__A2 (.I(_02641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06265__A2 (.I(_02641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06264__A2 (.I(_02641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06263__A2 (.I(_02641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06262__A2 (.I(_02641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06261__A2 (.I(_02641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06260__A2 (.I(_02641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06259__A2 (.I(_02641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06258__A2 (.I(_02641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06257__A2 (.I(_02641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06290__A2 (.I(_02651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06289__A2 (.I(_02651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06288__A2 (.I(_02651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06287__A2 (.I(_02651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06286__A2 (.I(_02651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06285__A2 (.I(_02651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06284__A2 (.I(_02651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06283__A2 (.I(_02651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06282__A2 (.I(_02651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06281__A2 (.I(_02651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06280__A2 (.I(_02651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06279__A2 (.I(_02651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06278__A2 (.I(_02651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06277__A2 (.I(_02651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06276__A2 (.I(_02651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06275__A2 (.I(_02651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08782__A2 (.I(_02660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08730__A1 (.I(_02660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07563__A1 (.I(_02660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07136__A2 (.I(_02660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07100__A1 (.I(_02660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06851__A1 (.I(_02660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06790__A2 (.I(_02660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06609__A2 (.I(_02660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06292__A2 (.I(_02660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06309__A2 (.I(_02662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06308__A2 (.I(_02662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06307__A2 (.I(_02662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06306__A2 (.I(_02662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06305__A2 (.I(_02662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06304__A2 (.I(_02662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06303__A2 (.I(_02662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06302__A2 (.I(_02662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06301__A2 (.I(_02662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06300__A2 (.I(_02662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06299__A2 (.I(_02662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06298__A2 (.I(_02662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06297__A2 (.I(_02662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06296__A2 (.I(_02662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06295__A2 (.I(_02662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06294__A2 (.I(_02662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09155__A1 (.I(_02671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08924__A2 (.I(_02671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07747__A2 (.I(_02671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07581__A1 (.I(_02671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07466__A2 (.I(_02671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07118__A1 (.I(_02671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06869__A1 (.I(_02671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06645__A2 (.I(_02671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06311__A2 (.I(_02671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06328__A2 (.I(_02673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06327__A2 (.I(_02673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06326__A2 (.I(_02673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06325__A2 (.I(_02673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06324__A2 (.I(_02673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06323__A2 (.I(_02673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06322__A2 (.I(_02673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06321__A2 (.I(_02673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06320__A2 (.I(_02673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06319__A2 (.I(_02673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06318__A2 (.I(_02673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06317__A2 (.I(_02673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06316__A2 (.I(_02673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06315__A2 (.I(_02673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06314__A2 (.I(_02673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06313__A2 (.I(_02673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09137__A2 (.I(_02682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09047__A1 (.I(_02682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08748__A2 (.I(_02682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07951__A1 (.I(_02682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07765__A2 (.I(_02682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07430__A1 (.I(_02682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06887__A2 (.I(_02682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06717__A2 (.I(_02682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06332__A1 (.I(_02682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09217__A1 (.I(_02684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07322__A2 (.I(_02684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07030__A2 (.I(_02684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07012__A2 (.I(_02684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06994__A1 (.I(_02684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06976__A2 (.I(_02684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06958__A1 (.I(_02684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06940__A1 (.I(_02684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06922__A2 (.I(_02684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06869__A2 (.I(_02684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06851__A2 (.I(_02684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06833__A2 (.I(_02684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06815__A1 (.I(_02684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06426__A2 (.I(_02684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06388__A2 (.I(_02684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06332__A2 (.I(_02684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06349__A2 (.I(_02686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06348__A2 (.I(_02686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06347__A2 (.I(_02686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06346__A2 (.I(_02686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06345__A2 (.I(_02686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06344__A2 (.I(_02686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06343__A2 (.I(_02686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06342__A2 (.I(_02686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06341__A2 (.I(_02686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06340__A2 (.I(_02686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06339__A2 (.I(_02686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06338__A2 (.I(_02686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06337__A2 (.I(_02686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06336__A2 (.I(_02686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06335__A2 (.I(_02686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06334__A2 (.I(_02686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09524__A2 (.I(_02695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09435__A2 (.I(_02695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09083__A1 (.I(_02695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07863__A1 (.I(_02695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07304__A1 (.I(_02695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07179__A2 (.I(_02695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07048__A2 (.I(_02695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06940__A2 (.I(_02695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06351__A2 (.I(_02695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06368__A2 (.I(_02697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06367__A2 (.I(_02697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06366__A2 (.I(_02697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06365__A2 (.I(_02697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06364__A2 (.I(_02697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06363__A2 (.I(_02697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06362__A2 (.I(_02697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06361__A2 (.I(_02697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06360__A2 (.I(_02697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06359__A2 (.I(_02697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06358__A2 (.I(_02697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06357__A2 (.I(_02697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06356__A2 (.I(_02697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06355__A2 (.I(_02697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06354__A2 (.I(_02697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06353__A2 (.I(_02697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09399__A2 (.I(_02706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09217__A2 (.I(_02706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09119__A1 (.I(_02706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07898__A2 (.I(_02706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07692__A2 (.I(_02706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07599__A1 (.I(_02706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06663__A2 (.I(_02706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06591__A1 (.I(_02706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06370__A2 (.I(_02706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06387__A2 (.I(_02708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06386__A2 (.I(_02708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06385__A2 (.I(_02708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06384__A2 (.I(_02708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06383__A2 (.I(_02708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06382__A2 (.I(_02708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06381__A2 (.I(_02708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06380__A2 (.I(_02708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06379__A2 (.I(_02708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06378__A2 (.I(_02708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06377__A2 (.I(_02708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06376__A2 (.I(_02708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06375__A2 (.I(_02708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06374__A2 (.I(_02708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06373__A2 (.I(_02708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06372__A2 (.I(_02708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06405__A2 (.I(_02718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06404__A2 (.I(_02718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06403__A2 (.I(_02718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06402__A2 (.I(_02718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06401__A2 (.I(_02718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06400__A2 (.I(_02718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06399__A2 (.I(_02718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06398__A2 (.I(_02718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06397__A2 (.I(_02718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06396__A2 (.I(_02718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06395__A2 (.I(_02718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06394__A2 (.I(_02718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06393__A2 (.I(_02718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06392__A2 (.I(_02718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06391__A2 (.I(_02718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06390__A2 (.I(_02718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09306__A1 (.I(_02727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09065__A2 (.I(_02727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08883__A2 (.I(_02727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08544__A2 (.I(_02727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07527__A1 (.I(_02727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07233__A1 (.I(_02727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07065__A2 (.I(_02727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06815__A2 (.I(_02727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06407__A2 (.I(_02727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06424__A2 (.I(_02729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06423__A2 (.I(_02729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06422__A2 (.I(_02729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06421__A2 (.I(_02729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06420__A2 (.I(_02729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06419__A2 (.I(_02729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06418__A2 (.I(_02729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06417__A2 (.I(_02729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06416__A2 (.I(_02729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06415__A2 (.I(_02729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06414__A2 (.I(_02729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06413__A2 (.I(_02729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06412__A2 (.I(_02729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06411__A2 (.I(_02729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06410__A2 (.I(_02729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06409__A2 (.I(_02729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06774__A1 (.I(_02738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06756__A1 (.I(_02738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06738__A1 (.I(_02738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06720__A1 (.I(_02738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06702__A1 (.I(_02738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06666__A1 (.I(_02738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06648__A1 (.I(_02738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06630__A1 (.I(_02738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06612__A1 (.I(_02738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06594__A1 (.I(_02738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06576__A1 (.I(_02738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06557__A1 (.I(_02738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06538__A1 (.I(_02738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06519__A1 (.I(_02738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06501__A1 (.I(_02738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06429__A1 (.I(_02738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06450__A2 (.I(_02740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06449__A2 (.I(_02740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06447__A2 (.I(_02740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06446__A2 (.I(_02740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06444__A2 (.I(_02740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06443__A2 (.I(_02740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06441__A2 (.I(_02740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06440__A2 (.I(_02740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06438__A2 (.I(_02740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06437__A2 (.I(_02740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06435__A2 (.I(_02740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06434__A2 (.I(_02740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06432__A2 (.I(_02740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06431__A2 (.I(_02740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06429__A2 (.I(_02740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06428__A2 (.I(_02740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06776__A1 (.I(_02742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06758__A1 (.I(_02742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06740__A1 (.I(_02742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06722__A1 (.I(_02742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06704__A1 (.I(_02742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06668__A1 (.I(_02742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06650__A1 (.I(_02742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06632__A1 (.I(_02742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06614__A1 (.I(_02742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06596__A1 (.I(_02742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06578__A1 (.I(_02742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06559__A1 (.I(_02742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06540__A1 (.I(_02742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06521__A1 (.I(_02742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06503__A1 (.I(_02742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06432__A1 (.I(_02742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06778__A1 (.I(_02744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06760__A1 (.I(_02744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06742__A1 (.I(_02744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06724__A1 (.I(_02744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06706__A1 (.I(_02744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06670__A1 (.I(_02744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06652__A1 (.I(_02744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06634__A1 (.I(_02744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06616__A1 (.I(_02744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06598__A1 (.I(_02744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06580__A1 (.I(_02744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06561__A1 (.I(_02744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06542__A1 (.I(_02744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06523__A1 (.I(_02744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06505__A1 (.I(_02744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06435__A1 (.I(_02744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06780__A1 (.I(_02746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06762__A1 (.I(_02746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06744__A1 (.I(_02746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06726__A1 (.I(_02746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06708__A1 (.I(_02746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06672__A1 (.I(_02746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06654__A1 (.I(_02746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06636__A1 (.I(_02746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06618__A1 (.I(_02746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06600__A1 (.I(_02746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06582__A1 (.I(_02746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06563__A1 (.I(_02746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06544__A1 (.I(_02746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06525__A1 (.I(_02746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06507__A1 (.I(_02746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06438__A1 (.I(_02746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06782__A1 (.I(_02748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06764__A1 (.I(_02748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06746__A1 (.I(_02748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06728__A1 (.I(_02748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06710__A1 (.I(_02748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06674__A1 (.I(_02748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06656__A1 (.I(_02748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06638__A1 (.I(_02748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06620__A1 (.I(_02748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06602__A1 (.I(_02748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06584__A1 (.I(_02748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06565__A1 (.I(_02748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06546__A1 (.I(_02748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06527__A1 (.I(_02748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06509__A1 (.I(_02748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06441__A1 (.I(_02748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06784__A1 (.I(_02750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06766__A1 (.I(_02750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06748__A1 (.I(_02750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06730__A1 (.I(_02750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06712__A1 (.I(_02750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06676__A1 (.I(_02750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06658__A1 (.I(_02750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06640__A1 (.I(_02750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06622__A1 (.I(_02750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06604__A1 (.I(_02750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06586__A1 (.I(_02750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06567__A1 (.I(_02750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06548__A1 (.I(_02750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06529__A1 (.I(_02750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06511__A1 (.I(_02750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06444__A1 (.I(_02750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06786__A1 (.I(_02752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06768__A1 (.I(_02752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06750__A1 (.I(_02752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06732__A1 (.I(_02752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06714__A1 (.I(_02752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06678__A1 (.I(_02752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06660__A1 (.I(_02752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06642__A1 (.I(_02752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06624__A1 (.I(_02752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06606__A1 (.I(_02752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06588__A1 (.I(_02752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06569__A1 (.I(_02752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06550__A1 (.I(_02752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06531__A1 (.I(_02752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06513__A1 (.I(_02752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06447__A1 (.I(_02752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06788__A1 (.I(_02754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06770__A1 (.I(_02754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06752__A1 (.I(_02754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06734__A1 (.I(_02754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06716__A1 (.I(_02754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06680__A1 (.I(_02754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06662__A1 (.I(_02754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06644__A1 (.I(_02754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06626__A1 (.I(_02754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06608__A1 (.I(_02754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06590__A1 (.I(_02754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06571__A1 (.I(_02754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06552__A1 (.I(_02754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06533__A1 (.I(_02754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06515__A1 (.I(_02754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06450__A1 (.I(_02754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06466__S (.I(_02756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06464__S (.I(_02756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06462__S (.I(_02756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06460__S (.I(_02756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06458__S (.I(_02756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06456__S (.I(_02756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06454__S (.I(_02756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06452__S (.I(_02756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08430__A1 (.I(_02765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08408__A1 (.I(_02765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08401__A1 (.I(_02765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08396__A1 (.I(_02765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08375__A1 (.I(_02765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08201__A1 (.I(_02765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08196__A1 (.I(_02765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08185__A1 (.I(_02765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08178__A1 (.I(_02765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08167__A1 (.I(_02765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08159__A1 (.I(_02765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08154__A1 (.I(_02765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08151__A1 (.I(_02765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08147__A1 (.I(_02765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06470__A1 (.I(_02765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08447__B (.I(_02767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06471__I (.I(_02767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08801__A1 (.I(_02768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08511__A1 (.I(_02768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08504__A2 (.I(_02768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08495__A2 (.I(_02768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08485__A2 (.I(_02768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08421__B2 (.I(_02768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08382__A1 (.I(_02768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08355__A2 (.I(_02768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08340__A1 (.I(_02768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08275__B2 (.I(_02768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08261__A1 (.I(_02768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08246__C (.I(_02768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08228__A2 (.I(_02768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08214__A1 (.I(_02768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08140__I (.I(_02768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06472__B (.I(_02768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09570__A1 (.I(_02769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06494__A1 (.I(_02769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06488__A1 (.I(_02769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06473__A2 (.I(_02769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06475__A2 (.I(_02770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08629__A2 (.I(_02773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08628__C (.I(_02773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08626__A2 (.I(_02773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07671__A2 (.I(_02773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06478__A2 (.I(_02773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08041__A2 (.I(_02774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08038__A1 (.I(_02774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08034__A2 (.I(_02774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08033__A1 (.I(_02774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08025__B (.I(_02774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08024__A2 (.I(_02774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08018__B (.I(_02774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08017__A2 (.I(_02774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08011__A2 (.I(_02774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08009__A2 (.I(_02774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06482__A1 (.I(_02774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08046__B2 (.I(_02779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06484__A3 (.I(_02779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08120__A2 (.I(_02781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08118__A2 (.I(_02781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08115__A2 (.I(_02781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08106__A2 (.I(_02781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08103__A1 (.I(_02781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08039__A1 (.I(_02781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08029__A2 (.I(_02781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08028__B (.I(_02781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08022__A2 (.I(_02781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08021__B (.I(_02781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08011__B (.I(_02781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06486__B (.I(_02781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09571__A1 (.I(_02783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07684__I (.I(_02783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06494__A2 (.I(_02783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06488__A2 (.I(_02783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06515__A2 (.I(_02791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06514__A2 (.I(_02791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06513__A2 (.I(_02791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06512__A2 (.I(_02791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06511__A2 (.I(_02791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06510__A2 (.I(_02791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06509__A2 (.I(_02791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06508__A2 (.I(_02791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06507__A2 (.I(_02791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06506__A2 (.I(_02791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06505__A2 (.I(_02791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06504__A2 (.I(_02791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06503__A2 (.I(_02791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06502__A2 (.I(_02791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06501__A2 (.I(_02791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06500__A2 (.I(_02791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06533__A2 (.I(_02801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06532__A2 (.I(_02801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06531__A2 (.I(_02801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06530__A2 (.I(_02801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06529__A2 (.I(_02801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06528__A2 (.I(_02801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06527__A2 (.I(_02801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06526__A2 (.I(_02801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06525__A2 (.I(_02801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06524__A2 (.I(_02801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06523__A2 (.I(_02801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06522__A2 (.I(_02801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06521__A2 (.I(_02801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06520__A2 (.I(_02801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06519__A2 (.I(_02801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06518__A2 (.I(_02801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09453__A2 (.I(_02810_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09342__A2 (.I(_02810_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09029__A1 (.I(_02810_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07881__A2 (.I(_02810_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07820__A1 (.I(_02810_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07340__A1 (.I(_02810_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07154__A2 (.I(_02810_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06958__A2 (.I(_02810_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06535__A2 (.I(_02810_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06552__A2 (.I(_02812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06551__A2 (.I(_02812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06550__A2 (.I(_02812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06549__A2 (.I(_02812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06548__A2 (.I(_02812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06547__A2 (.I(_02812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06546__A2 (.I(_02812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06545__A2 (.I(_02812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06544__A2 (.I(_02812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06543__A2 (.I(_02812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06542__A2 (.I(_02812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06541__A2 (.I(_02812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06540__A2 (.I(_02812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06539__A2 (.I(_02812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06538__A2 (.I(_02812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06537__A2 (.I(_02812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08289__A2 (.I(_02821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08122__A2 (.I(_02821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07969__A2 (.I(_02821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07951__A2 (.I(_02821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07933__A2 (.I(_02821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07915__A2 (.I(_02821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07863__A2 (.I(_02821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07845__A1 (.I(_02821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07820__A2 (.I(_02821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07801__A2 (.I(_02821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07599__A2 (.I(_02821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07581__A2 (.I(_02821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07563__A2 (.I(_02821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07545__A2 (.I(_02821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07527__A2 (.I(_02821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06554__A2 (.I(_02821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06571__A2 (.I(_02823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06570__A2 (.I(_02823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06569__A2 (.I(_02823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06568__A2 (.I(_02823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06567__A2 (.I(_02823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06566__A2 (.I(_02823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06565__A2 (.I(_02823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06564__A2 (.I(_02823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06563__A2 (.I(_02823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06562__A2 (.I(_02823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06561__A2 (.I(_02823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06560__A2 (.I(_02823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06559__A2 (.I(_02823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06558__A2 (.I(_02823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06557__A2 (.I(_02823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06556__A2 (.I(_02823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07509__A2 (.I(_02832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07448__A2 (.I(_02832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07430__A2 (.I(_02832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07412__A2 (.I(_02832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07394__A2 (.I(_02832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07376__A1 (.I(_02832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07358__A2 (.I(_02832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07340__A2 (.I(_02832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07304__A2 (.I(_02832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07268__A2 (.I(_02832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07233__A2 (.I(_02832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07118__A2 (.I(_02832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07100__A2 (.I(_02832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07082__A2 (.I(_02832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06591__A2 (.I(_02832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06573__A2 (.I(_02832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06590__A2 (.I(_02834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06589__A2 (.I(_02834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06588__A2 (.I(_02834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06587__A2 (.I(_02834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06586__A2 (.I(_02834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06585__A2 (.I(_02834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06584__A2 (.I(_02834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06583__A2 (.I(_02834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06582__A2 (.I(_02834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06581__A2 (.I(_02834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06580__A2 (.I(_02834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06579__A2 (.I(_02834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06578__A2 (.I(_02834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06577__A2 (.I(_02834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06576__A2 (.I(_02834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06575__A2 (.I(_02834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06608__A2 (.I(_02844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06607__A2 (.I(_02844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06606__A2 (.I(_02844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06605__A2 (.I(_02844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06604__A2 (.I(_02844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06603__A2 (.I(_02844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06602__A2 (.I(_02844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06601__A2 (.I(_02844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06600__A2 (.I(_02844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06599__A2 (.I(_02844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06598__A2 (.I(_02844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06597__A2 (.I(_02844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06596__A2 (.I(_02844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06595__A2 (.I(_02844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06594__A2 (.I(_02844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06593__A2 (.I(_02844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06626__A2 (.I(_02854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06625__A2 (.I(_02854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06624__A2 (.I(_02854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06623__A2 (.I(_02854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06622__A2 (.I(_02854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06621__A2 (.I(_02854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06620__A2 (.I(_02854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06619__A2 (.I(_02854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06618__A2 (.I(_02854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06617__A2 (.I(_02854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06616__A2 (.I(_02854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06615__A2 (.I(_02854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06614__A2 (.I(_02854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06613__A2 (.I(_02854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06612__A2 (.I(_02854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06611__A2 (.I(_02854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06644__A2 (.I(_02864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06643__A2 (.I(_02864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06642__A2 (.I(_02864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06641__A2 (.I(_02864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06640__A2 (.I(_02864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06639__A2 (.I(_02864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06638__A2 (.I(_02864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06637__A2 (.I(_02864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06636__A2 (.I(_02864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06635__A2 (.I(_02864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06634__A2 (.I(_02864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06633__A2 (.I(_02864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06632__A2 (.I(_02864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06631__A2 (.I(_02864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06630__A2 (.I(_02864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06629__A2 (.I(_02864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06662__A2 (.I(_02874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06661__A2 (.I(_02874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06660__A2 (.I(_02874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06659__A2 (.I(_02874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06658__A2 (.I(_02874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06657__A2 (.I(_02874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06656__A2 (.I(_02874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06655__A2 (.I(_02874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06654__A2 (.I(_02874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06653__A2 (.I(_02874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06652__A2 (.I(_02874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06651__A2 (.I(_02874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06650__A2 (.I(_02874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06649__A2 (.I(_02874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06648__A2 (.I(_02874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06647__A2 (.I(_02874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06680__A2 (.I(_02884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06679__A2 (.I(_02884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06678__A2 (.I(_02884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06677__A2 (.I(_02884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06676__A2 (.I(_02884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06675__A2 (.I(_02884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06674__A2 (.I(_02884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06673__A2 (.I(_02884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06672__A2 (.I(_02884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06671__A2 (.I(_02884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06670__A2 (.I(_02884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06669__A2 (.I(_02884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06668__A2 (.I(_02884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06667__A2 (.I(_02884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06666__A2 (.I(_02884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06665__A2 (.I(_02884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09288__A2 (.I(_02893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08993__A1 (.I(_02893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07845__A2 (.I(_02893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07617__A2 (.I(_02893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07484__A2 (.I(_02893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07376__A2 (.I(_02893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07215__A2 (.I(_02893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06994__A2 (.I(_02893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06682__A2 (.I(_02893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06697__S (.I(_02894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06695__S (.I(_02894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06693__S (.I(_02894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06691__S (.I(_02894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06689__S (.I(_02894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06687__S (.I(_02894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06685__S (.I(_02894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06683__S (.I(_02894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06716__A2 (.I(_02904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06715__A2 (.I(_02904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06714__A2 (.I(_02904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06713__A2 (.I(_02904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06712__A2 (.I(_02904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06711__A2 (.I(_02904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06710__A2 (.I(_02904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06709__A2 (.I(_02904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06708__A2 (.I(_02904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06707__A2 (.I(_02904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06706__A2 (.I(_02904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06705__A2 (.I(_02904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06704__A2 (.I(_02904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06703__A2 (.I(_02904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06702__A2 (.I(_02904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06701__A2 (.I(_02904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06734__A2 (.I(_02914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06733__A2 (.I(_02914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06732__A2 (.I(_02914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06731__A2 (.I(_02914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06730__A2 (.I(_02914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06729__A2 (.I(_02914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06728__A2 (.I(_02914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06727__A2 (.I(_02914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06726__A2 (.I(_02914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06725__A2 (.I(_02914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06724__A2 (.I(_02914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06723__A2 (.I(_02914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06722__A2 (.I(_02914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06721__A2 (.I(_02914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06720__A2 (.I(_02914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06719__A2 (.I(_02914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06752__A2 (.I(_02924_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06751__A2 (.I(_02924_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06750__A2 (.I(_02924_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06749__A2 (.I(_02924_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06748__A2 (.I(_02924_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06747__A2 (.I(_02924_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06746__A2 (.I(_02924_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06745__A2 (.I(_02924_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06744__A2 (.I(_02924_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06743__A2 (.I(_02924_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06742__A2 (.I(_02924_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06741__A2 (.I(_02924_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06740__A2 (.I(_02924_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06739__A2 (.I(_02924_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06738__A2 (.I(_02924_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06737__A2 (.I(_02924_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06770__A2 (.I(_02934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06769__A2 (.I(_02934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06768__A2 (.I(_02934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06767__A2 (.I(_02934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06766__A2 (.I(_02934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06765__A2 (.I(_02934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06764__A2 (.I(_02934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06763__A2 (.I(_02934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06762__A2 (.I(_02934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06761__A2 (.I(_02934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06760__A2 (.I(_02934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06759__A2 (.I(_02934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06758__A2 (.I(_02934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06757__A2 (.I(_02934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06756__A2 (.I(_02934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06755__A2 (.I(_02934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06788__A2 (.I(_02944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06787__A2 (.I(_02944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06786__A2 (.I(_02944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06785__A2 (.I(_02944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06784__A2 (.I(_02944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06783__A2 (.I(_02944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06782__A2 (.I(_02944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06781__A2 (.I(_02944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06780__A2 (.I(_02944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06779__A2 (.I(_02944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06778__A2 (.I(_02944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06777__A2 (.I(_02944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06776__A2 (.I(_02944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06775__A2 (.I(_02944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06774__A2 (.I(_02944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06773__A2 (.I(_02944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07121__A1 (.I(_02953_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07103__A1 (.I(_02953_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07085__A1 (.I(_02953_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07033__A1 (.I(_02953_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07015__A1 (.I(_02953_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06997__A1 (.I(_02953_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06979__A1 (.I(_02953_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06961__A1 (.I(_02953_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06943__A1 (.I(_02953_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06925__A1 (.I(_02953_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06890__A1 (.I(_02953_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06872__A1 (.I(_02953_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06854__A1 (.I(_02953_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06836__A1 (.I(_02953_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06818__A1 (.I(_02953_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06793__A1 (.I(_02953_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06814__A2 (.I(_02955_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06813__A2 (.I(_02955_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06811__A2 (.I(_02955_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06810__A2 (.I(_02955_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06808__A2 (.I(_02955_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06807__A2 (.I(_02955_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06805__A2 (.I(_02955_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06804__A2 (.I(_02955_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06802__A2 (.I(_02955_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06801__A2 (.I(_02955_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06799__A2 (.I(_02955_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06798__A2 (.I(_02955_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06796__A2 (.I(_02955_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06795__A2 (.I(_02955_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06793__A2 (.I(_02955_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06792__A2 (.I(_02955_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07123__A1 (.I(_02957_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07105__A1 (.I(_02957_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07087__A1 (.I(_02957_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07035__A1 (.I(_02957_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07017__A1 (.I(_02957_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06999__A1 (.I(_02957_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06981__A1 (.I(_02957_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06963__A1 (.I(_02957_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06945__A1 (.I(_02957_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06927__A1 (.I(_02957_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06892__A1 (.I(_02957_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06874__A1 (.I(_02957_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06856__A1 (.I(_02957_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06838__A1 (.I(_02957_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06820__A1 (.I(_02957_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06796__A1 (.I(_02957_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07125__A1 (.I(_02959_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07107__A1 (.I(_02959_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07089__A1 (.I(_02959_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07037__A1 (.I(_02959_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07019__A1 (.I(_02959_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07001__A1 (.I(_02959_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06983__A1 (.I(_02959_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06965__A1 (.I(_02959_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06947__A1 (.I(_02959_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06929__A1 (.I(_02959_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06894__A1 (.I(_02959_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06876__A1 (.I(_02959_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06858__A1 (.I(_02959_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06840__A1 (.I(_02959_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06822__A1 (.I(_02959_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06799__A1 (.I(_02959_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07127__A1 (.I(_02961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07109__A1 (.I(_02961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07091__A1 (.I(_02961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07039__A1 (.I(_02961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07021__A1 (.I(_02961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07003__A1 (.I(_02961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06985__A1 (.I(_02961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06967__A1 (.I(_02961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06949__A1 (.I(_02961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06931__A1 (.I(_02961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06896__A1 (.I(_02961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06878__A1 (.I(_02961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06860__A1 (.I(_02961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06842__A1 (.I(_02961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06824__A1 (.I(_02961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06802__A1 (.I(_02961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07129__A1 (.I(_02963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07111__A1 (.I(_02963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07093__A1 (.I(_02963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07041__A1 (.I(_02963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07023__A1 (.I(_02963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07005__A1 (.I(_02963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06987__A1 (.I(_02963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06969__A1 (.I(_02963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06951__A1 (.I(_02963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06933__A1 (.I(_02963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06898__A1 (.I(_02963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06880__A1 (.I(_02963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06862__A1 (.I(_02963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06844__A1 (.I(_02963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06826__A1 (.I(_02963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06805__A1 (.I(_02963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07131__A1 (.I(_02965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07113__A1 (.I(_02965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07095__A1 (.I(_02965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07043__A1 (.I(_02965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07025__A1 (.I(_02965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07007__A1 (.I(_02965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06989__A1 (.I(_02965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06971__A1 (.I(_02965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06953__A1 (.I(_02965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06935__A1 (.I(_02965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06900__A1 (.I(_02965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06882__A1 (.I(_02965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06864__A1 (.I(_02965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06846__A1 (.I(_02965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06828__A1 (.I(_02965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06808__A1 (.I(_02965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07133__A1 (.I(_02967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07115__A1 (.I(_02967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07097__A1 (.I(_02967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07045__A1 (.I(_02967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07027__A1 (.I(_02967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07009__A1 (.I(_02967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06991__A1 (.I(_02967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06973__A1 (.I(_02967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06955__A1 (.I(_02967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06937__A1 (.I(_02967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06902__A1 (.I(_02967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06884__A1 (.I(_02967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06866__A1 (.I(_02967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06848__A1 (.I(_02967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06830__A1 (.I(_02967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06811__A1 (.I(_02967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07135__A1 (.I(_02969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07117__A1 (.I(_02969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07099__A1 (.I(_02969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07047__A1 (.I(_02969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07029__A1 (.I(_02969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07011__A1 (.I(_02969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06993__A1 (.I(_02969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06975__A1 (.I(_02969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06957__A1 (.I(_02969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06939__A1 (.I(_02969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06904__A1 (.I(_02969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06886__A1 (.I(_02969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06868__A1 (.I(_02969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06850__A1 (.I(_02969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06832__A1 (.I(_02969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06814__A1 (.I(_02969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06832__A2 (.I(_02972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06831__A2 (.I(_02972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06830__A2 (.I(_02972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06829__A2 (.I(_02972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06828__A2 (.I(_02972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06827__A2 (.I(_02972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06826__A2 (.I(_02972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06825__A2 (.I(_02972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06824__A2 (.I(_02972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06823__A2 (.I(_02972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06822__A2 (.I(_02972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06821__A2 (.I(_02972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06820__A2 (.I(_02972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06819__A2 (.I(_02972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06818__A2 (.I(_02972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06817__A2 (.I(_02972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06850__A2 (.I(_02982_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06849__A2 (.I(_02982_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06848__A2 (.I(_02982_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06847__A2 (.I(_02982_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06846__A2 (.I(_02982_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06845__A2 (.I(_02982_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06844__A2 (.I(_02982_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06843__A2 (.I(_02982_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06842__A2 (.I(_02982_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06841__A2 (.I(_02982_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06840__A2 (.I(_02982_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06839__A2 (.I(_02982_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06838__A2 (.I(_02982_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06837__A2 (.I(_02982_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06836__A2 (.I(_02982_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06835__A2 (.I(_02982_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06868__A2 (.I(_02992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06867__A2 (.I(_02992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06866__A2 (.I(_02992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06865__A2 (.I(_02992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06864__A2 (.I(_02992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06863__A2 (.I(_02992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06862__A2 (.I(_02992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06861__A2 (.I(_02992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06860__A2 (.I(_02992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06859__A2 (.I(_02992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06858__A2 (.I(_02992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06857__A2 (.I(_02992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06856__A2 (.I(_02992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06855__A2 (.I(_02992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06854__A2 (.I(_02992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06853__A2 (.I(_02992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06886__A2 (.I(_03002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06885__A2 (.I(_03002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06884__A2 (.I(_03002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06883__A2 (.I(_03002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06882__A2 (.I(_03002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06881__A2 (.I(_03002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06880__A2 (.I(_03002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06879__A2 (.I(_03002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06878__A2 (.I(_03002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06877__A2 (.I(_03002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06876__A2 (.I(_03002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06875__A2 (.I(_03002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06874__A2 (.I(_03002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06873__A2 (.I(_03002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06872__A2 (.I(_03002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06871__A2 (.I(_03002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06904__A2 (.I(_03012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06903__A2 (.I(_03012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06902__A2 (.I(_03012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06901__A2 (.I(_03012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06900__A2 (.I(_03012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06899__A2 (.I(_03012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06898__A2 (.I(_03012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06897__A2 (.I(_03012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06896__A2 (.I(_03012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06895__A2 (.I(_03012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06894__A2 (.I(_03012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06893__A2 (.I(_03012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06892__A2 (.I(_03012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06891__A2 (.I(_03012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06890__A2 (.I(_03012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06889__A2 (.I(_03012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06920__S (.I(_03021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06918__S (.I(_03021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06916__S (.I(_03021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06914__S (.I(_03021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06912__S (.I(_03021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06910__S (.I(_03021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06908__S (.I(_03021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06906__S (.I(_03021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06939__A2 (.I(_03031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06938__A2 (.I(_03031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06937__A2 (.I(_03031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06936__A2 (.I(_03031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06935__A2 (.I(_03031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06934__A2 (.I(_03031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06933__A2 (.I(_03031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06932__A2 (.I(_03031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06931__A2 (.I(_03031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06930__A2 (.I(_03031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06929__A2 (.I(_03031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06928__A2 (.I(_03031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06927__A2 (.I(_03031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06926__A2 (.I(_03031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06925__A2 (.I(_03031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06924__A2 (.I(_03031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06957__A2 (.I(_03041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06956__A2 (.I(_03041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06955__A2 (.I(_03041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06954__A2 (.I(_03041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06953__A2 (.I(_03041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06952__A2 (.I(_03041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06951__A2 (.I(_03041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06950__A2 (.I(_03041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06949__A2 (.I(_03041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06948__A2 (.I(_03041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06947__A2 (.I(_03041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06946__A2 (.I(_03041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06945__A2 (.I(_03041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06944__A2 (.I(_03041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06943__A2 (.I(_03041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06942__A2 (.I(_03041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06975__A2 (.I(_03051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06974__A2 (.I(_03051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06973__A2 (.I(_03051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06972__A2 (.I(_03051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06971__A2 (.I(_03051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06970__A2 (.I(_03051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06969__A2 (.I(_03051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06968__A2 (.I(_03051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06967__A2 (.I(_03051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06966__A2 (.I(_03051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06965__A2 (.I(_03051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06964__A2 (.I(_03051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06963__A2 (.I(_03051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06962__A2 (.I(_03051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06961__A2 (.I(_03051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06960__A2 (.I(_03051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06993__A2 (.I(_03061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06992__A2 (.I(_03061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06991__A2 (.I(_03061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06990__A2 (.I(_03061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06989__A2 (.I(_03061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06988__A2 (.I(_03061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06987__A2 (.I(_03061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06986__A2 (.I(_03061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06985__A2 (.I(_03061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06984__A2 (.I(_03061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06983__A2 (.I(_03061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06982__A2 (.I(_03061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06981__A2 (.I(_03061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06980__A2 (.I(_03061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06979__A2 (.I(_03061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06978__A2 (.I(_03061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07011__A2 (.I(_03071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07010__A2 (.I(_03071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07009__A2 (.I(_03071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07008__A2 (.I(_03071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07007__A2 (.I(_03071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07006__A2 (.I(_03071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07005__A2 (.I(_03071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07004__A2 (.I(_03071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07003__A2 (.I(_03071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07002__A2 (.I(_03071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07001__A2 (.I(_03071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07000__A2 (.I(_03071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06999__A2 (.I(_03071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06998__A2 (.I(_03071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06997__A2 (.I(_03071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06996__A2 (.I(_03071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07029__A2 (.I(_03081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07028__A2 (.I(_03081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07027__A2 (.I(_03081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07026__A2 (.I(_03081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07025__A2 (.I(_03081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07024__A2 (.I(_03081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07023__A2 (.I(_03081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07022__A2 (.I(_03081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07021__A2 (.I(_03081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07020__A2 (.I(_03081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07019__A2 (.I(_03081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07018__A2 (.I(_03081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07017__A2 (.I(_03081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07016__A2 (.I(_03081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07015__A2 (.I(_03081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07014__A2 (.I(_03081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07047__A2 (.I(_03091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07046__A2 (.I(_03091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07045__A2 (.I(_03091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07044__A2 (.I(_03091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07043__A2 (.I(_03091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07042__A2 (.I(_03091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07041__A2 (.I(_03091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07040__A2 (.I(_03091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07039__A2 (.I(_03091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07038__A2 (.I(_03091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07037__A2 (.I(_03091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07036__A2 (.I(_03091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07035__A2 (.I(_03091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07034__A2 (.I(_03091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07033__A2 (.I(_03091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07032__A2 (.I(_03091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07063__S (.I(_03100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07061__S (.I(_03100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07059__S (.I(_03100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07057__S (.I(_03100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07055__S (.I(_03100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07053__S (.I(_03100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07051__S (.I(_03100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07049__S (.I(_03100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07080__S (.I(_03109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07078__S (.I(_03109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07076__S (.I(_03109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07074__S (.I(_03109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07072__S (.I(_03109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07070__S (.I(_03109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07068__S (.I(_03109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07066__S (.I(_03109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07099__A2 (.I(_03119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07098__A2 (.I(_03119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07097__A2 (.I(_03119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07096__A2 (.I(_03119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07095__A2 (.I(_03119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07094__A2 (.I(_03119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07093__A2 (.I(_03119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07092__A2 (.I(_03119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07091__A2 (.I(_03119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07090__A2 (.I(_03119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07089__A2 (.I(_03119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07088__A2 (.I(_03119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07087__A2 (.I(_03119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07086__A2 (.I(_03119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07085__A2 (.I(_03119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07084__A2 (.I(_03119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07117__A2 (.I(_03129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07116__A2 (.I(_03129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07115__A2 (.I(_03129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07114__A2 (.I(_03129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07113__A2 (.I(_03129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07112__A2 (.I(_03129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07111__A2 (.I(_03129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07110__A2 (.I(_03129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07109__A2 (.I(_03129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07108__A2 (.I(_03129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07107__A2 (.I(_03129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07106__A2 (.I(_03129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07105__A2 (.I(_03129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07104__A2 (.I(_03129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07103__A2 (.I(_03129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07102__A2 (.I(_03129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07135__A2 (.I(_03139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07134__A2 (.I(_03139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07133__A2 (.I(_03139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07132__A2 (.I(_03139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07131__A2 (.I(_03139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07130__A2 (.I(_03139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07129__A2 (.I(_03139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07128__A2 (.I(_03139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07127__A2 (.I(_03139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07126__A2 (.I(_03139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07125__A2 (.I(_03139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07124__A2 (.I(_03139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07123__A2 (.I(_03139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07122__A2 (.I(_03139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07121__A2 (.I(_03139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07120__A2 (.I(_03139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07151__S (.I(_03148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07149__S (.I(_03148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07147__S (.I(_03148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07145__S (.I(_03148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07143__S (.I(_03148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07141__S (.I(_03148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07139__S (.I(_03148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07137__S (.I(_03148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07451__A1 (.I(_03157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07433__A1 (.I(_03157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07415__A1 (.I(_03157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07397__A1 (.I(_03157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07379__A1 (.I(_03157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07361__A1 (.I(_03157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07343__A1 (.I(_03157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07325__A1 (.I(_03157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07307__A1 (.I(_03157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07289__A1 (.I(_03157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07271__A1 (.I(_03157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07236__A1 (.I(_03157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07218__A1 (.I(_03157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07200__A1 (.I(_03157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07182__A1 (.I(_03157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07157__A1 (.I(_03157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07178__A2 (.I(_03159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07177__A2 (.I(_03159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07175__A2 (.I(_03159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07174__A2 (.I(_03159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07172__A2 (.I(_03159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07171__A2 (.I(_03159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07169__A2 (.I(_03159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07168__A2 (.I(_03159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07166__A2 (.I(_03159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07165__A2 (.I(_03159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07163__A2 (.I(_03159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07162__A2 (.I(_03159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07160__A2 (.I(_03159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07159__A2 (.I(_03159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07157__A2 (.I(_03159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07156__A2 (.I(_03159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07453__A1 (.I(_03161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07435__A1 (.I(_03161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07417__A1 (.I(_03161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07399__A1 (.I(_03161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07381__A1 (.I(_03161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07363__A1 (.I(_03161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07345__A1 (.I(_03161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07327__A1 (.I(_03161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07309__A1 (.I(_03161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07291__A1 (.I(_03161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07273__A1 (.I(_03161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07238__A1 (.I(_03161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07220__A1 (.I(_03161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07202__A1 (.I(_03161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07184__A1 (.I(_03161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07160__A1 (.I(_03161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07455__A1 (.I(_03163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07437__A1 (.I(_03163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07419__A1 (.I(_03163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07401__A1 (.I(_03163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07383__A1 (.I(_03163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07365__A1 (.I(_03163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07347__A1 (.I(_03163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07329__A1 (.I(_03163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07311__A1 (.I(_03163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07293__A1 (.I(_03163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07275__A1 (.I(_03163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07240__A1 (.I(_03163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07222__A1 (.I(_03163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07204__A1 (.I(_03163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07186__A1 (.I(_03163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07163__A1 (.I(_03163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07457__A1 (.I(_03165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07439__A1 (.I(_03165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07421__A1 (.I(_03165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07403__A1 (.I(_03165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07385__A1 (.I(_03165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07367__A1 (.I(_03165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07349__A1 (.I(_03165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07331__A1 (.I(_03165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07313__A1 (.I(_03165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07295__A1 (.I(_03165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07277__A1 (.I(_03165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07242__A1 (.I(_03165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07224__A1 (.I(_03165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07206__A1 (.I(_03165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07188__A1 (.I(_03165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07166__A1 (.I(_03165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07459__A1 (.I(_03167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07441__A1 (.I(_03167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07423__A1 (.I(_03167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07405__A1 (.I(_03167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07387__A1 (.I(_03167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07369__A1 (.I(_03167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07351__A1 (.I(_03167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07333__A1 (.I(_03167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07315__A1 (.I(_03167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07297__A1 (.I(_03167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07279__A1 (.I(_03167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07244__A1 (.I(_03167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07226__A1 (.I(_03167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07208__A1 (.I(_03167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07190__A1 (.I(_03167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07169__A1 (.I(_03167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07461__A1 (.I(_03169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07443__A1 (.I(_03169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07425__A1 (.I(_03169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07407__A1 (.I(_03169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07389__A1 (.I(_03169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07371__A1 (.I(_03169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07353__A1 (.I(_03169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07335__A1 (.I(_03169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07317__A1 (.I(_03169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07299__A1 (.I(_03169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07281__A1 (.I(_03169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07246__A1 (.I(_03169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07228__A1 (.I(_03169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07210__A1 (.I(_03169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07192__A1 (.I(_03169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07172__A1 (.I(_03169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07463__A1 (.I(_03171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07445__A1 (.I(_03171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07427__A1 (.I(_03171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07409__A1 (.I(_03171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07391__A1 (.I(_03171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07373__A1 (.I(_03171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07355__A1 (.I(_03171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07337__A1 (.I(_03171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07319__A1 (.I(_03171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07301__A1 (.I(_03171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07283__A1 (.I(_03171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07248__A1 (.I(_03171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07230__A1 (.I(_03171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07212__A1 (.I(_03171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07194__A1 (.I(_03171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07175__A1 (.I(_03171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07465__A1 (.I(_03173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07447__A1 (.I(_03173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07429__A1 (.I(_03173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07411__A1 (.I(_03173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07393__A1 (.I(_03173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07375__A1 (.I(_03173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07357__A1 (.I(_03173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07339__A1 (.I(_03173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07321__A1 (.I(_03173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07303__A1 (.I(_03173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07285__A1 (.I(_03173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07250__A1 (.I(_03173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07232__A1 (.I(_03173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07214__A1 (.I(_03173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07196__A1 (.I(_03173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07178__A1 (.I(_03173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07196__A2 (.I(_03176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07195__A2 (.I(_03176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07194__A2 (.I(_03176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07193__A2 (.I(_03176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07192__A2 (.I(_03176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07191__A2 (.I(_03176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07190__A2 (.I(_03176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07189__A2 (.I(_03176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07188__A2 (.I(_03176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07187__A2 (.I(_03176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07186__A2 (.I(_03176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07185__A2 (.I(_03176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07184__A2 (.I(_03176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07183__A2 (.I(_03176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07182__A2 (.I(_03176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07181__A2 (.I(_03176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07214__A2 (.I(_03186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07213__A2 (.I(_03186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07212__A2 (.I(_03186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07211__A2 (.I(_03186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07210__A2 (.I(_03186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07209__A2 (.I(_03186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07208__A2 (.I(_03186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07207__A2 (.I(_03186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07206__A2 (.I(_03186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07205__A2 (.I(_03186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07204__A2 (.I(_03186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07203__A2 (.I(_03186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07202__A2 (.I(_03186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07201__A2 (.I(_03186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07200__A2 (.I(_03186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07199__A2 (.I(_03186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07232__A2 (.I(_03196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07231__A2 (.I(_03196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07230__A2 (.I(_03196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07229__A2 (.I(_03196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07228__A2 (.I(_03196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07227__A2 (.I(_03196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07226__A2 (.I(_03196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07225__A2 (.I(_03196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07224__A2 (.I(_03196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07223__A2 (.I(_03196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07222__A2 (.I(_03196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07221__A2 (.I(_03196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07220__A2 (.I(_03196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07219__A2 (.I(_03196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07218__A2 (.I(_03196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07217__A2 (.I(_03196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07250__A2 (.I(_03206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07249__A2 (.I(_03206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07248__A2 (.I(_03206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07247__A2 (.I(_03206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07246__A2 (.I(_03206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07245__A2 (.I(_03206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07244__A2 (.I(_03206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07243__A2 (.I(_03206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07242__A2 (.I(_03206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07241__A2 (.I(_03206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07240__A2 (.I(_03206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07239__A2 (.I(_03206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07238__A2 (.I(_03206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07237__A2 (.I(_03206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07236__A2 (.I(_03206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07235__A2 (.I(_03206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07266__S (.I(_03215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07264__S (.I(_03215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07262__S (.I(_03215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07260__S (.I(_03215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07258__S (.I(_03215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07256__S (.I(_03215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07254__S (.I(_03215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07252__S (.I(_03215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07285__A2 (.I(_03225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07284__A2 (.I(_03225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07283__A2 (.I(_03225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07282__A2 (.I(_03225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07281__A2 (.I(_03225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07280__A2 (.I(_03225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07279__A2 (.I(_03225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07278__A2 (.I(_03225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07277__A2 (.I(_03225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07276__A2 (.I(_03225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07275__A2 (.I(_03225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07274__A2 (.I(_03225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07273__A2 (.I(_03225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07272__A2 (.I(_03225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07271__A2 (.I(_03225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07270__A2 (.I(_03225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07303__A2 (.I(_03235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07302__A2 (.I(_03235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07301__A2 (.I(_03235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07300__A2 (.I(_03235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07299__A2 (.I(_03235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07298__A2 (.I(_03235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07297__A2 (.I(_03235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07296__A2 (.I(_03235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07295__A2 (.I(_03235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07294__A2 (.I(_03235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07293__A2 (.I(_03235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07292__A2 (.I(_03235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07291__A2 (.I(_03235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07290__A2 (.I(_03235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07289__A2 (.I(_03235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07288__A2 (.I(_03235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07321__A2 (.I(_03245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07320__A2 (.I(_03245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07319__A2 (.I(_03245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07318__A2 (.I(_03245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07317__A2 (.I(_03245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07316__A2 (.I(_03245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07315__A2 (.I(_03245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07314__A2 (.I(_03245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07313__A2 (.I(_03245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07312__A2 (.I(_03245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07311__A2 (.I(_03245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07310__A2 (.I(_03245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07309__A2 (.I(_03245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07308__A2 (.I(_03245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07307__A2 (.I(_03245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07306__A2 (.I(_03245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07339__A2 (.I(_03255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07338__A2 (.I(_03255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07337__A2 (.I(_03255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07336__A2 (.I(_03255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07335__A2 (.I(_03255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07334__A2 (.I(_03255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07333__A2 (.I(_03255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07332__A2 (.I(_03255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07331__A2 (.I(_03255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07330__A2 (.I(_03255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07329__A2 (.I(_03255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07328__A2 (.I(_03255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07327__A2 (.I(_03255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07326__A2 (.I(_03255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07325__A2 (.I(_03255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07324__A2 (.I(_03255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07357__A2 (.I(_03265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07356__A2 (.I(_03265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07355__A2 (.I(_03265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07354__A2 (.I(_03265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07353__A2 (.I(_03265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07352__A2 (.I(_03265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07351__A2 (.I(_03265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07350__A2 (.I(_03265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07349__A2 (.I(_03265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07348__A2 (.I(_03265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07347__A2 (.I(_03265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07346__A2 (.I(_03265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07345__A2 (.I(_03265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07344__A2 (.I(_03265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07343__A2 (.I(_03265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07342__A2 (.I(_03265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07375__A2 (.I(_03275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07374__A2 (.I(_03275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07373__A2 (.I(_03275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07372__A2 (.I(_03275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07371__A2 (.I(_03275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07370__A2 (.I(_03275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07369__A2 (.I(_03275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07368__A2 (.I(_03275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07367__A2 (.I(_03275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07366__A2 (.I(_03275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07365__A2 (.I(_03275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07364__A2 (.I(_03275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07363__A2 (.I(_03275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07362__A2 (.I(_03275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07361__A2 (.I(_03275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07360__A2 (.I(_03275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07393__A2 (.I(_03285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07392__A2 (.I(_03285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07391__A2 (.I(_03285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07390__A2 (.I(_03285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07389__A2 (.I(_03285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07388__A2 (.I(_03285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07387__A2 (.I(_03285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07386__A2 (.I(_03285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07385__A2 (.I(_03285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07384__A2 (.I(_03285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07383__A2 (.I(_03285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07382__A2 (.I(_03285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07381__A2 (.I(_03285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07380__A2 (.I(_03285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07379__A2 (.I(_03285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07378__A2 (.I(_03285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07411__A2 (.I(_03295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07410__A2 (.I(_03295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07409__A2 (.I(_03295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07408__A2 (.I(_03295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07407__A2 (.I(_03295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07406__A2 (.I(_03295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07405__A2 (.I(_03295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07404__A2 (.I(_03295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07403__A2 (.I(_03295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07402__A2 (.I(_03295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07401__A2 (.I(_03295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07400__A2 (.I(_03295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07399__A2 (.I(_03295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07398__A2 (.I(_03295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07397__A2 (.I(_03295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07396__A2 (.I(_03295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07429__A2 (.I(_03305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07428__A2 (.I(_03305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07427__A2 (.I(_03305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07426__A2 (.I(_03305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07425__A2 (.I(_03305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07424__A2 (.I(_03305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07423__A2 (.I(_03305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07422__A2 (.I(_03305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07421__A2 (.I(_03305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07420__A2 (.I(_03305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07419__A2 (.I(_03305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07418__A2 (.I(_03305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07417__A2 (.I(_03305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07416__A2 (.I(_03305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07415__A2 (.I(_03305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07414__A2 (.I(_03305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07447__A2 (.I(_03315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07446__A2 (.I(_03315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07445__A2 (.I(_03315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07444__A2 (.I(_03315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07443__A2 (.I(_03315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07442__A2 (.I(_03315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07441__A2 (.I(_03315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07440__A2 (.I(_03315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07439__A2 (.I(_03315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07438__A2 (.I(_03315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07437__A2 (.I(_03315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07436__A2 (.I(_03315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07435__A2 (.I(_03315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07434__A2 (.I(_03315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07433__A2 (.I(_03315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07432__A2 (.I(_03315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07465__A2 (.I(_03325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07464__A2 (.I(_03325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07463__A2 (.I(_03325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07462__A2 (.I(_03325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07461__A2 (.I(_03325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07460__A2 (.I(_03325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07459__A2 (.I(_03325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07458__A2 (.I(_03325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07457__A2 (.I(_03325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07456__A2 (.I(_03325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07455__A2 (.I(_03325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07454__A2 (.I(_03325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07453__A2 (.I(_03325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07452__A2 (.I(_03325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07451__A2 (.I(_03325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07450__A2 (.I(_03325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07481__S (.I(_03334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07479__S (.I(_03334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07477__S (.I(_03334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07475__S (.I(_03334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07473__S (.I(_03334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07471__S (.I(_03334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07469__S (.I(_03334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07467__S (.I(_03334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07804__A1 (.I(_03343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07786__A1 (.I(_03343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07768__A1 (.I(_03343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07750__A1 (.I(_03343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07713__A1 (.I(_03343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07695__A1 (.I(_03343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07656__A1 (.I(_03343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07638__A1 (.I(_03343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07620__A1 (.I(_03343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07602__A1 (.I(_03343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07584__A1 (.I(_03343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07566__A1 (.I(_03343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07548__A1 (.I(_03343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07530__A1 (.I(_03343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07512__A1 (.I(_03343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07487__A1 (.I(_03343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07508__A2 (.I(_03345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07507__A2 (.I(_03345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07505__A2 (.I(_03345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07504__A2 (.I(_03345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07502__A2 (.I(_03345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07501__A2 (.I(_03345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07499__A2 (.I(_03345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07498__A2 (.I(_03345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07496__A2 (.I(_03345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07495__A2 (.I(_03345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07493__A2 (.I(_03345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07492__A2 (.I(_03345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07490__A2 (.I(_03345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07489__A2 (.I(_03345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07487__A2 (.I(_03345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07486__A2 (.I(_03345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07806__A1 (.I(_03347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07788__A1 (.I(_03347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07770__A1 (.I(_03347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07752__A1 (.I(_03347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07715__A1 (.I(_03347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07697__A1 (.I(_03347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07658__A1 (.I(_03347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07640__A1 (.I(_03347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07622__A1 (.I(_03347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07604__A1 (.I(_03347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07586__A1 (.I(_03347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07568__A1 (.I(_03347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07550__A1 (.I(_03347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07532__A1 (.I(_03347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07514__A1 (.I(_03347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07490__A1 (.I(_03347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07808__A1 (.I(_03349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07790__A1 (.I(_03349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07772__A1 (.I(_03349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07754__A1 (.I(_03349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07717__A1 (.I(_03349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07699__A1 (.I(_03349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07660__A1 (.I(_03349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07642__A1 (.I(_03349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07624__A1 (.I(_03349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07606__A1 (.I(_03349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07588__A1 (.I(_03349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07570__A1 (.I(_03349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07552__A1 (.I(_03349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07534__A1 (.I(_03349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07516__A1 (.I(_03349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07493__A1 (.I(_03349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07810__A1 (.I(_03351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07792__A1 (.I(_03351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07774__A1 (.I(_03351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07756__A1 (.I(_03351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07719__A1 (.I(_03351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07701__A1 (.I(_03351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07662__A1 (.I(_03351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07644__A1 (.I(_03351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07626__A1 (.I(_03351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07608__A1 (.I(_03351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07590__A1 (.I(_03351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07572__A1 (.I(_03351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07554__A1 (.I(_03351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07536__A1 (.I(_03351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07518__A1 (.I(_03351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07496__A1 (.I(_03351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07812__A1 (.I(_03353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07794__A1 (.I(_03353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07776__A1 (.I(_03353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07758__A1 (.I(_03353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07721__A1 (.I(_03353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07703__A1 (.I(_03353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07664__A1 (.I(_03353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07646__A1 (.I(_03353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07628__A1 (.I(_03353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07610__A1 (.I(_03353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07592__A1 (.I(_03353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07574__A1 (.I(_03353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07556__A1 (.I(_03353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07538__A1 (.I(_03353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07520__A1 (.I(_03353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07499__A1 (.I(_03353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07814__A1 (.I(_03355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07796__A1 (.I(_03355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07778__A1 (.I(_03355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07760__A1 (.I(_03355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07723__A1 (.I(_03355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07705__A1 (.I(_03355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07666__A1 (.I(_03355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07648__A1 (.I(_03355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07630__A1 (.I(_03355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07612__A1 (.I(_03355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07594__A1 (.I(_03355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07576__A1 (.I(_03355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07558__A1 (.I(_03355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07540__A1 (.I(_03355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07522__A1 (.I(_03355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07502__A1 (.I(_03355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07816__A1 (.I(_03357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07798__A1 (.I(_03357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07780__A1 (.I(_03357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07762__A1 (.I(_03357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07725__A1 (.I(_03357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07707__A1 (.I(_03357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07668__A1 (.I(_03357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07650__A1 (.I(_03357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07632__A1 (.I(_03357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07614__A1 (.I(_03357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07596__A1 (.I(_03357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07578__A1 (.I(_03357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07560__A1 (.I(_03357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07542__A1 (.I(_03357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07524__A1 (.I(_03357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07505__A1 (.I(_03357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07818__A1 (.I(_03359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07800__A1 (.I(_03359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07782__A1 (.I(_03359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07764__A1 (.I(_03359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07727__A1 (.I(_03359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07709__A1 (.I(_03359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07670__A1 (.I(_03359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07652__A1 (.I(_03359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07634__A1 (.I(_03359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07616__A1 (.I(_03359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07598__A1 (.I(_03359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07580__A1 (.I(_03359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07562__A1 (.I(_03359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07544__A1 (.I(_03359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07526__A1 (.I(_03359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07508__A1 (.I(_03359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07526__A2 (.I(_03362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07525__A2 (.I(_03362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07524__A2 (.I(_03362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07523__A2 (.I(_03362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07522__A2 (.I(_03362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07521__A2 (.I(_03362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07520__A2 (.I(_03362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07519__A2 (.I(_03362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07518__A2 (.I(_03362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07517__A2 (.I(_03362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07516__A2 (.I(_03362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07515__A2 (.I(_03362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07514__A2 (.I(_03362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07513__A2 (.I(_03362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07512__A2 (.I(_03362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07511__A2 (.I(_03362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07544__A2 (.I(_03372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07543__A2 (.I(_03372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07542__A2 (.I(_03372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07541__A2 (.I(_03372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07540__A2 (.I(_03372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07539__A2 (.I(_03372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07538__A2 (.I(_03372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07537__A2 (.I(_03372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07536__A2 (.I(_03372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07535__A2 (.I(_03372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07534__A2 (.I(_03372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07533__A2 (.I(_03372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07532__A2 (.I(_03372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07531__A2 (.I(_03372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07530__A2 (.I(_03372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07529__A2 (.I(_03372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07562__A2 (.I(_03382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07561__A2 (.I(_03382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07560__A2 (.I(_03382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07559__A2 (.I(_03382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07558__A2 (.I(_03382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07557__A2 (.I(_03382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07556__A2 (.I(_03382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07555__A2 (.I(_03382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07554__A2 (.I(_03382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07553__A2 (.I(_03382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07552__A2 (.I(_03382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07551__A2 (.I(_03382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07550__A2 (.I(_03382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07549__A2 (.I(_03382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07548__A2 (.I(_03382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07547__A2 (.I(_03382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07580__A2 (.I(_03392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07579__A2 (.I(_03392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07578__A2 (.I(_03392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07577__A2 (.I(_03392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07576__A2 (.I(_03392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07575__A2 (.I(_03392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07574__A2 (.I(_03392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07573__A2 (.I(_03392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07572__A2 (.I(_03392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07571__A2 (.I(_03392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07570__A2 (.I(_03392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07569__A2 (.I(_03392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07568__A2 (.I(_03392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07567__A2 (.I(_03392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07566__A2 (.I(_03392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07565__A2 (.I(_03392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07598__A2 (.I(_03402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07597__A2 (.I(_03402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07596__A2 (.I(_03402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07595__A2 (.I(_03402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07594__A2 (.I(_03402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07593__A2 (.I(_03402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07592__A2 (.I(_03402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07591__A2 (.I(_03402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07590__A2 (.I(_03402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07589__A2 (.I(_03402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07588__A2 (.I(_03402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07587__A2 (.I(_03402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07586__A2 (.I(_03402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07585__A2 (.I(_03402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07584__A2 (.I(_03402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07583__A2 (.I(_03402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07616__A2 (.I(_03412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07615__A2 (.I(_03412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07614__A2 (.I(_03412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07613__A2 (.I(_03412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07612__A2 (.I(_03412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07611__A2 (.I(_03412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07610__A2 (.I(_03412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07609__A2 (.I(_03412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07608__A2 (.I(_03412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07607__A2 (.I(_03412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07606__A2 (.I(_03412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07605__A2 (.I(_03412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07604__A2 (.I(_03412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07603__A2 (.I(_03412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07602__A2 (.I(_03412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07601__A2 (.I(_03412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07634__A2 (.I(_03422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07633__A2 (.I(_03422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07632__A2 (.I(_03422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07631__A2 (.I(_03422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07630__A2 (.I(_03422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07629__A2 (.I(_03422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07628__A2 (.I(_03422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07627__A2 (.I(_03422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07626__A2 (.I(_03422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07625__A2 (.I(_03422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07624__A2 (.I(_03422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07623__A2 (.I(_03422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07622__A2 (.I(_03422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07621__A2 (.I(_03422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07620__A2 (.I(_03422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07619__A2 (.I(_03422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07652__A2 (.I(_03432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07651__A2 (.I(_03432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07650__A2 (.I(_03432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07649__A2 (.I(_03432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07648__A2 (.I(_03432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07647__A2 (.I(_03432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07646__A2 (.I(_03432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07645__A2 (.I(_03432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07644__A2 (.I(_03432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07643__A2 (.I(_03432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07642__A2 (.I(_03432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07641__A2 (.I(_03432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07640__A2 (.I(_03432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07639__A2 (.I(_03432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07638__A2 (.I(_03432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07637__A2 (.I(_03432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07670__A2 (.I(_03442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07669__A2 (.I(_03442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07668__A2 (.I(_03442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07667__A2 (.I(_03442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07666__A2 (.I(_03442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07665__A2 (.I(_03442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07664__A2 (.I(_03442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07663__A2 (.I(_03442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07662__A2 (.I(_03442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07661__A2 (.I(_03442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07660__A2 (.I(_03442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07659__A2 (.I(_03442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07658__A2 (.I(_03442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07657__A2 (.I(_03442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07656__A2 (.I(_03442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07655__A2 (.I(_03442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09387__A2 (.I(_03454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07679__A2 (.I(_03454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07678__A2 (.I(_03454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07677__A2 (.I(_03454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07676__A3 (.I(_03454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09560__A2 (.I(_03458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09397__A2 (.I(_03458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07745__A2 (.I(_03458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07731__A2 (.I(_03458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07729__A2 (.I(_03458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07683__A2 (.I(_03458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07709__A2 (.I(_03465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07708__A2 (.I(_03465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07707__A2 (.I(_03465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07706__A2 (.I(_03465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07705__A2 (.I(_03465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07704__A2 (.I(_03465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07703__A2 (.I(_03465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07702__A2 (.I(_03465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07701__A2 (.I(_03465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07700__A2 (.I(_03465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07699__A2 (.I(_03465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07698__A2 (.I(_03465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07697__A2 (.I(_03465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07696__A2 (.I(_03465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07695__A2 (.I(_03465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07694__A2 (.I(_03465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07727__A2 (.I(_03475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07726__A2 (.I(_03475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07725__A2 (.I(_03475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07724__A2 (.I(_03475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07723__A2 (.I(_03475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07722__A2 (.I(_03475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07721__A2 (.I(_03475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07720__A2 (.I(_03475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07719__A2 (.I(_03475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07718__A2 (.I(_03475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07717__A2 (.I(_03475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07716__A2 (.I(_03475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07715__A2 (.I(_03475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07714__A2 (.I(_03475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07713__A2 (.I(_03475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07712__A2 (.I(_03475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07764__A2 (.I(_03500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07763__A2 (.I(_03500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07762__A2 (.I(_03500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07761__A2 (.I(_03500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07760__A2 (.I(_03500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07759__A2 (.I(_03500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07758__A2 (.I(_03500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07757__A2 (.I(_03500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07756__A2 (.I(_03500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07755__A2 (.I(_03500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07754__A2 (.I(_03500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07753__A2 (.I(_03500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07752__A2 (.I(_03500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07751__A2 (.I(_03500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07750__A2 (.I(_03500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07749__A2 (.I(_03500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07782__A2 (.I(_03510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07781__A2 (.I(_03510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07780__A2 (.I(_03510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07779__A2 (.I(_03510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07778__A2 (.I(_03510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07777__A2 (.I(_03510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07776__A2 (.I(_03510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07775__A2 (.I(_03510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07774__A2 (.I(_03510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07773__A2 (.I(_03510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07772__A2 (.I(_03510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07771__A2 (.I(_03510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07770__A2 (.I(_03510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07769__A2 (.I(_03510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07768__A2 (.I(_03510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07767__A2 (.I(_03510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07800__A2 (.I(_03520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07799__A2 (.I(_03520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07798__A2 (.I(_03520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07797__A2 (.I(_03520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07796__A2 (.I(_03520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07795__A2 (.I(_03520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07794__A2 (.I(_03520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07793__A2 (.I(_03520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07792__A2 (.I(_03520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07791__A2 (.I(_03520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07790__A2 (.I(_03520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07789__A2 (.I(_03520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07788__A2 (.I(_03520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07787__A2 (.I(_03520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07786__A2 (.I(_03520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07785__A2 (.I(_03520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07818__A2 (.I(_03530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07817__A2 (.I(_03530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07816__A2 (.I(_03530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07815__A2 (.I(_03530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07814__A2 (.I(_03530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07813__A2 (.I(_03530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07812__A2 (.I(_03530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07811__A2 (.I(_03530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07810__A2 (.I(_03530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07809__A2 (.I(_03530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07808__A2 (.I(_03530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07807__A2 (.I(_03530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07806__A2 (.I(_03530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07805__A2 (.I(_03530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07804__A2 (.I(_03530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07803__A2 (.I(_03530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08842__A1 (.I(_03539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08785__A1 (.I(_03539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08733__A1 (.I(_03539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08639__A1 (.I(_03539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08547__A1 (.I(_03539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08529__A1 (.I(_03539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08292__A1 (.I(_03539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08125__A1 (.I(_03539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07990__A1 (.I(_03539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07972__A1 (.I(_03539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07954__A1 (.I(_03539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07936__A1 (.I(_03539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07918__A1 (.I(_03539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07866__A1 (.I(_03539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07848__A1 (.I(_03539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07823__A1 (.I(_03539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07844__A2 (.I(_03541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07843__A2 (.I(_03541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07841__A2 (.I(_03541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07840__A2 (.I(_03541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07838__A2 (.I(_03541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07837__A2 (.I(_03541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07835__A2 (.I(_03541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07834__A2 (.I(_03541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07832__A2 (.I(_03541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07831__A2 (.I(_03541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07829__A2 (.I(_03541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07828__A2 (.I(_03541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07826__A2 (.I(_03541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07825__A2 (.I(_03541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07823__A2 (.I(_03541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07822__A2 (.I(_03541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08844__A1 (.I(_03543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08787__A1 (.I(_03543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08735__A1 (.I(_03543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08641__A1 (.I(_03543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08549__A1 (.I(_03543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08531__A1 (.I(_03543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08294__A1 (.I(_03543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08127__A1 (.I(_03543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07992__A1 (.I(_03543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07974__A1 (.I(_03543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07956__A1 (.I(_03543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07938__A1 (.I(_03543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07920__A1 (.I(_03543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07868__A1 (.I(_03543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07850__A1 (.I(_03543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07826__A1 (.I(_03543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08846__A1 (.I(_03545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08789__A1 (.I(_03545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08737__A1 (.I(_03545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08643__A1 (.I(_03545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08551__A1 (.I(_03545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08533__A1 (.I(_03545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08296__A1 (.I(_03545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08129__A1 (.I(_03545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07994__A1 (.I(_03545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07976__A1 (.I(_03545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07958__A1 (.I(_03545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07940__A1 (.I(_03545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07922__A1 (.I(_03545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07870__A1 (.I(_03545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07852__A1 (.I(_03545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07829__A1 (.I(_03545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08848__A1 (.I(_03547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08791__A1 (.I(_03547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08739__A1 (.I(_03547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08645__A1 (.I(_03547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08553__A1 (.I(_03547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08535__A1 (.I(_03547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08298__A1 (.I(_03547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08131__A1 (.I(_03547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07996__A1 (.I(_03547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07978__A1 (.I(_03547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07960__A1 (.I(_03547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07942__A1 (.I(_03547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07924__A1 (.I(_03547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07872__A1 (.I(_03547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07854__A1 (.I(_03547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07832__A1 (.I(_03547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08850__A1 (.I(_03549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08793__A1 (.I(_03549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08741__A1 (.I(_03549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08647__A1 (.I(_03549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08555__A1 (.I(_03549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08537__A1 (.I(_03549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08300__A1 (.I(_03549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08133__A1 (.I(_03549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07998__A1 (.I(_03549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07980__A1 (.I(_03549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07962__A1 (.I(_03549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07944__A1 (.I(_03549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07926__A1 (.I(_03549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07874__A1 (.I(_03549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07856__A1 (.I(_03549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07835__A1 (.I(_03549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08852__A1 (.I(_03551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08795__A1 (.I(_03551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08743__A1 (.I(_03551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08649__A1 (.I(_03551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08557__A1 (.I(_03551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08539__A1 (.I(_03551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08302__A1 (.I(_03551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08135__A1 (.I(_03551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08000__A1 (.I(_03551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07982__A1 (.I(_03551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07964__A1 (.I(_03551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07946__A1 (.I(_03551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07928__A1 (.I(_03551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07876__A1 (.I(_03551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07858__A1 (.I(_03551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07838__A1 (.I(_03551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08854__A1 (.I(_03553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08797__A1 (.I(_03553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08745__A1 (.I(_03553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08651__A1 (.I(_03553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08559__A1 (.I(_03553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08541__A1 (.I(_03553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08304__A1 (.I(_03553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08137__A1 (.I(_03553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08002__A1 (.I(_03553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07984__A1 (.I(_03553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07966__A1 (.I(_03553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07948__A1 (.I(_03553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07930__A1 (.I(_03553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07878__A1 (.I(_03553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07860__A1 (.I(_03553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07841__A1 (.I(_03553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08856__A1 (.I(_03555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08799__A1 (.I(_03555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08747__A1 (.I(_03555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08653__A1 (.I(_03555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08561__A1 (.I(_03555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08543__A1 (.I(_03555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08306__A1 (.I(_03555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08139__A1 (.I(_03555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08004__A1 (.I(_03555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07986__A1 (.I(_03555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07968__A1 (.I(_03555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07950__A1 (.I(_03555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07932__A1 (.I(_03555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07880__A1 (.I(_03555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07862__A1 (.I(_03555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07844__A1 (.I(_03555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07862__A2 (.I(_03558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07861__A2 (.I(_03558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07860__A2 (.I(_03558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07859__A2 (.I(_03558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07858__A2 (.I(_03558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07857__A2 (.I(_03558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07856__A2 (.I(_03558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07855__A2 (.I(_03558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07854__A2 (.I(_03558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07853__A2 (.I(_03558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07852__A2 (.I(_03558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07851__A2 (.I(_03558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07850__A2 (.I(_03558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07849__A2 (.I(_03558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07848__A2 (.I(_03558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07847__A2 (.I(_03558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07880__A2 (.I(_03568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07879__A2 (.I(_03568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07878__A2 (.I(_03568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07877__A2 (.I(_03568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07876__A2 (.I(_03568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07875__A2 (.I(_03568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07874__A2 (.I(_03568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07873__A2 (.I(_03568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07872__A2 (.I(_03568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07871__A2 (.I(_03568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07870__A2 (.I(_03568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07869__A2 (.I(_03568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07868__A2 (.I(_03568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07867__A2 (.I(_03568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07866__A2 (.I(_03568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07865__A2 (.I(_03568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07896__S (.I(_03577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07894__S (.I(_03577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07892__S (.I(_03577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07890__S (.I(_03577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07888__S (.I(_03577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07886__S (.I(_03577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07884__S (.I(_03577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07882__S (.I(_03577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07913__S (.I(_03586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07911__S (.I(_03586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07909__S (.I(_03586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07907__S (.I(_03586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07905__S (.I(_03586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07903__S (.I(_03586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07901__S (.I(_03586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07899__S (.I(_03586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07932__A2 (.I(_03596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07931__A2 (.I(_03596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07930__A2 (.I(_03596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07929__A2 (.I(_03596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07928__A2 (.I(_03596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07927__A2 (.I(_03596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07926__A2 (.I(_03596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07925__A2 (.I(_03596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07924__A2 (.I(_03596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07923__A2 (.I(_03596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07922__A2 (.I(_03596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07921__A2 (.I(_03596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07920__A2 (.I(_03596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07919__A2 (.I(_03596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07918__A2 (.I(_03596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07917__A2 (.I(_03596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07950__A2 (.I(_03606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07949__A2 (.I(_03606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07948__A2 (.I(_03606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07947__A2 (.I(_03606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07946__A2 (.I(_03606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07945__A2 (.I(_03606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07944__A2 (.I(_03606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07943__A2 (.I(_03606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07942__A2 (.I(_03606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07941__A2 (.I(_03606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07940__A2 (.I(_03606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07939__A2 (.I(_03606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07938__A2 (.I(_03606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07937__A2 (.I(_03606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07936__A2 (.I(_03606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07935__A2 (.I(_03606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07968__A2 (.I(_03616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07967__A2 (.I(_03616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07966__A2 (.I(_03616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07965__A2 (.I(_03616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07964__A2 (.I(_03616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07963__A2 (.I(_03616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07962__A2 (.I(_03616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07961__A2 (.I(_03616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07960__A2 (.I(_03616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07959__A2 (.I(_03616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07958__A2 (.I(_03616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07957__A2 (.I(_03616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07956__A2 (.I(_03616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07955__A2 (.I(_03616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07954__A2 (.I(_03616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07953__A2 (.I(_03616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07986__A2 (.I(_03626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07985__A2 (.I(_03626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07984__A2 (.I(_03626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07983__A2 (.I(_03626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07982__A2 (.I(_03626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07981__A2 (.I(_03626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07980__A2 (.I(_03626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07979__A2 (.I(_03626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07978__A2 (.I(_03626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07977__A2 (.I(_03626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07976__A2 (.I(_03626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07975__A2 (.I(_03626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07974__A2 (.I(_03626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07973__A2 (.I(_03626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07972__A2 (.I(_03626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07971__A2 (.I(_03626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08004__A2 (.I(_03636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08003__A2 (.I(_03636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08002__A2 (.I(_03636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08001__A2 (.I(_03636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08000__A2 (.I(_03636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07999__A2 (.I(_03636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07998__A2 (.I(_03636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07997__A2 (.I(_03636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07996__A2 (.I(_03636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07995__A2 (.I(_03636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07994__A2 (.I(_03636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07993__A2 (.I(_03636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07992__A2 (.I(_03636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07991__A2 (.I(_03636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07990__A2 (.I(_03636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07989__A2 (.I(_03636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08103__A2 (.I(_03648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08039__A2 (.I(_03648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08034__B (.I(_03648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08026__A1 (.I(_03648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08019__A1 (.I(_03648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08014__A2 (.I(_03648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08010__A1 (.I(_03648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08112__A2 (.I(_03653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08109__A2 (.I(_03653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08104__A2 (.I(_03653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08097__A2 (.I(_03653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08094__A2 (.I(_03653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08091__A2 (.I(_03653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08080__A2 (.I(_03653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08072__A2 (.I(_03653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08048__A2 (.I(_03653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08035__B (.I(_03653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08032__I (.I(_03653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08015__A2 (.I(_03653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08014__A1 (.I(_03653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08112__B1 (.I(_03654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08109__B1 (.I(_03654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08104__B1 (.I(_03654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08100__A2 (.I(_03654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08097__B1 (.I(_03654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08094__B1 (.I(_03654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08091__B1 (.I(_03654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08089__B1 (.I(_03654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08080__B1 (.I(_03654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08072__B1 (.I(_03654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08048__B1 (.I(_03654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08046__A2 (.I(_03654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08042__I (.I(_03654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08015__B1 (.I(_03654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08509__A2 (.I(_03668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08161__A2 (.I(_03668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08036__A1 (.I(_03668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08099__A2 (.I(_03669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08089__A2 (.I(_03669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08086__A2 (.I(_03669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08083__A2 (.I(_03669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08078__A2 (.I(_03669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08075__A2 (.I(_03669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08070__A2 (.I(_03669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08067__A2 (.I(_03669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08064__A2 (.I(_03669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08061__A2 (.I(_03669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08058__A2 (.I(_03669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08055__A2 (.I(_03669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08052__A2 (.I(_03669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08045__A2 (.I(_03669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08043__A2 (.I(_03669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08036__A2 (.I(_03669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08108__A2 (.I(_03676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08100__B1 (.I(_03676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08091__C1 (.I(_03676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08080__C1 (.I(_03676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08072__C1 (.I(_03676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08050__I (.I(_03676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08048__C1 (.I(_03676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08046__B1 (.I(_03676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08041__C (.I(_03676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08121__A2 (.I(_03678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08119__A2 (.I(_03678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08116__A2 (.I(_03678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08107__A2 (.I(_03678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08086__B1 (.I(_03678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08083__B1 (.I(_03678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08078__B1 (.I(_03678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08075__B1 (.I(_03678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08070__B1 (.I(_03678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08067__B1 (.I(_03678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08064__B1 (.I(_03678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08061__B1 (.I(_03678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08058__B1 (.I(_03678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08055__B1 (.I(_03678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08052__B1 (.I(_03678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08043__B1 (.I(_03678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08119__B1 (.I(_03683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08116__B1 (.I(_03683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08096__A2 (.I(_03683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08093__A2 (.I(_03683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08088__A2 (.I(_03683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08085__A2 (.I(_03683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08082__A2 (.I(_03683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08077__A2 (.I(_03683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08074__A2 (.I(_03683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08069__A2 (.I(_03683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08066__A2 (.I(_03683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08063__A2 (.I(_03683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08060__A2 (.I(_03683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08057__A2 (.I(_03683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08054__A2 (.I(_03683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08051__A2 (.I(_03683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08120__B1 (.I(_03718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08113__A2 (.I(_03718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08106__B1 (.I(_03718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08105__A2 (.I(_03718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08139__A2 (.I(_03731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08138__A2 (.I(_03731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08137__A2 (.I(_03731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08136__A2 (.I(_03731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08135__A2 (.I(_03731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08134__A2 (.I(_03731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08133__A2 (.I(_03731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08132__A2 (.I(_03731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08131__A2 (.I(_03731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08130__A2 (.I(_03731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08129__A2 (.I(_03731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08128__A2 (.I(_03731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08127__A2 (.I(_03731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08126__A2 (.I(_03731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08125__A2 (.I(_03731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08124__A2 (.I(_03731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08836__A1 (.I(_03740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08824__B2 (.I(_03740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08810__A1 (.I(_03740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08471__C (.I(_03740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08378__A2 (.I(_03740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08333__A2 (.I(_03740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08288__A2 (.I(_03740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08276__A2 (.I(_03740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08264__A2 (.I(_03740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08253__A2 (.I(_03740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08252__A1 (.I(_03740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08247__A2 (.I(_03740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08240__A2 (.I(_03740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08239__A1 (.I(_03740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08195__A2 (.I(_03740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08194__A1 (.I(_03740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08836__A2 (.I(_03741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08512__A1 (.I(_03741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08507__A1 (.I(_03741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08417__A1 (.I(_03741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08416__B (.I(_03741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08360__A1 (.I(_03741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08358__A1 (.I(_03741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08320__A1 (.I(_03741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08242__A1 (.I(_03741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08222__A1 (.I(_03741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08145__A1 (.I(_03741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08827__B2 (.I(_03742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08501__A1 (.I(_03742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08499__A1 (.I(_03742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08417__A2 (.I(_03742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08416__A1 (.I(_03742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08410__A1 (.I(_03742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08350__A1 (.I(_03742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08321__A1 (.I(_03742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08243__A1 (.I(_03742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08222__A2 (.I(_03742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08145__A2 (.I(_03742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08816__A1 (.I(_03743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08489__A1 (.I(_03743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08398__A1 (.I(_03743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08145__A3 (.I(_03743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08441__A1 (.I(_03744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08439__B2 (.I(_03744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08436__A1 (.I(_03744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08329__C2 (.I(_03744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08327__B2 (.I(_03744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08324__A1 (.I(_03744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08145__A4 (.I(_03744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08807__A1 (.I(_03747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08481__A1 (.I(_03747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08477__A1 (.I(_03747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08148__A2 (.I(_03747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08462__A1 (.I(_03751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08416__A2 (.I(_03751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08241__A1 (.I(_03751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08152__A2 (.I(_03751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08255__A1 (.I(_03752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08210__A1 (.I(_03752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08193__A1 (.I(_03752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08438__A1 (.I(_03754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08259__A1 (.I(_03754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08230__A1 (.I(_03754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08225__A1 (.I(_03754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08191__A1 (.I(_03754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08171__A1 (.I(_03754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08826__A1 (.I(_03755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08433__C (.I(_03755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08361__A1 (.I(_03755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08272__B2 (.I(_03755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08230__A2 (.I(_03755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08191__A2 (.I(_03755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08180__A2 (.I(_03755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08174__A2 (.I(_03755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08171__A2 (.I(_03755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08478__A1 (.I(_03756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08388__A1 (.I(_03756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08358__B2 (.I(_03756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08284__A1 (.I(_03756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08157__I (.I(_03756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08815__B2 (.I(_03757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08361__A2 (.I(_03757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08248__A1 (.I(_03757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08243__A2 (.I(_03757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08232__A1 (.I(_03757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08229__B2 (.I(_03757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08165__A1 (.I(_03757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08348__B (.I(_03759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08248__A2 (.I(_03759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08232__A2 (.I(_03759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08225__B2 (.I(_03759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08165__A2 (.I(_03759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08808__A1 (.I(_03761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08389__A1 (.I(_03761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08386__A1 (.I(_03761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08273__B2 (.I(_03761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08266__A1 (.I(_03761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08244__A1 (.I(_03761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08206__A1 (.I(_03761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08164__A1 (.I(_03761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08814__A1 (.I(_03762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08397__A1 (.I(_03762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08283__A1 (.I(_03762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08282__A1 (.I(_03762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08250__A1 (.I(_03762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08219__B1 (.I(_03762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08164__A2 (.I(_03762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08439__A1 (.I(_03763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08367__B (.I(_03763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08327__A1 (.I(_03763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08260__A1 (.I(_03763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08256__A1 (.I(_03763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08255__B2 (.I(_03763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08234__A1 (.I(_03763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08183__A1 (.I(_03763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08164__A3 (.I(_03763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08462__A2 (.I(_03765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08209__A1 (.I(_03765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08170__A1 (.I(_03765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08365__A2 (.I(_03767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08329__A1 (.I(_03767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08271__A1 (.I(_03767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08269__A1 (.I(_03767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08251__A1 (.I(_03767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08245__A2 (.I(_03767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08233__A1 (.I(_03767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08231__A1 (.I(_03767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08216__A2 (.I(_03767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08204__A1 (.I(_03767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08169__A1 (.I(_03767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08471__A1 (.I(_03768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08462__A3 (.I(_03768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08350__A2 (.I(_03768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08315__A2 (.I(_03768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08270__A1 (.I(_03768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08269__A2 (.I(_03768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08211__A2 (.I(_03768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08169__A2 (.I(_03768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08815__A2 (.I(_03769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08329__B1 (.I(_03769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08221__A1 (.I(_03769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08170__A2 (.I(_03769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08821__A2 (.I(_03770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08432__A3 (.I(_03770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08255__A2 (.I(_03770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08171__A3 (.I(_03770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08833__A1 (.I(_03773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08387__A1 (.I(_03773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08370__A2 (.I(_03773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08369__A1 (.I(_03773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08365__A1 (.I(_03773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08328__A1 (.I(_03773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08272__A1 (.I(_03773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08268__A1 (.I(_03773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08258__A1 (.I(_03773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08245__A1 (.I(_03773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08216__A1 (.I(_03773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08215__A1 (.I(_03773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08202__A1 (.I(_03773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08180__A1 (.I(_03773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08174__A1 (.I(_03773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08471__A2 (.I(_03774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08261__A2 (.I(_03774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08251__A2 (.I(_03774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08213__A1 (.I(_03774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08182__A1 (.I(_03774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08489__A2 (.I(_03776_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08476__A2 (.I(_03776_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08463__A2 (.I(_03776_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08435__A2 (.I(_03776_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08409__A1 (.I(_03776_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08351__A1 (.I(_03776_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08317__A2 (.I(_03776_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08315__A1 (.I(_03776_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08211__A1 (.I(_03776_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08187__A1 (.I(_03776_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08186__A1 (.I(_03776_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08179__A1 (.I(_03776_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08827__A1 (.I(_03778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08814__A2 (.I(_03778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08808__A2 (.I(_03778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08461__A1 (.I(_03778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08439__A2 (.I(_03778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08436__B2 (.I(_03778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08360__A2 (.I(_03778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08284__A2 (.I(_03778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08233__A2 (.I(_03778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08231__A2 (.I(_03778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08225__A2 (.I(_03778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08209__A2 (.I(_03778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08187__A2 (.I(_03778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08179__A2 (.I(_03778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08808__B1 (.I(_03779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08489__B1 (.I(_03779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08475__A1 (.I(_03779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08439__B1 (.I(_03779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08391__B2 (.I(_03779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08360__B1 (.I(_03779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08319__A1 (.I(_03779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08284__B1 (.I(_03779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08181__A1 (.I(_03779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08827__A2 (.I(_03780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08818__A1 (.I(_03780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08809__A1 (.I(_03780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08806__B (.I(_03780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08499__B (.I(_03780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08361__B1 (.I(_03780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08330__A1 (.I(_03780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08274__A1 (.I(_03780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08181__A2 (.I(_03780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08822__A1 (.I(_03782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08807__B2 (.I(_03782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08510__B (.I(_03782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08503__A1 (.I(_03782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08494__A1 (.I(_03782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08490__A1 (.I(_03782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08484__A1 (.I(_03782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08483__B (.I(_03782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08469__C (.I(_03782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08354__A1 (.I(_03782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08353__C (.I(_03782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08286__A2 (.I(_03782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08237__A1 (.I(_03782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08225__B1 (.I(_03782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08206__A2 (.I(_03782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08183__A2 (.I(_03782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08366__A1 (.I(_03785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08319__A2 (.I(_03785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08316__A1 (.I(_03785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08311__A1 (.I(_03785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08256__A2 (.I(_03785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08190__A1 (.I(_03785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08186__A2 (.I(_03785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08826__A2 (.I(_03786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08500__A1 (.I(_03786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08461__A2 (.I(_03786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08419__A2 (.I(_03786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08410__A2 (.I(_03786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08398__A2 (.I(_03786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08358__A2 (.I(_03786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08324__A2 (.I(_03786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08257__A1 (.I(_03786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08192__A1 (.I(_03786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08812__A1 (.I(_03788_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08808__B2 (.I(_03788_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08804__B (.I(_03788_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08479__B (.I(_03788_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08476__A1 (.I(_03788_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08419__A1 (.I(_03788_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08391__A1 (.I(_03788_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08389__B2 (.I(_03788_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08310__A2 (.I(_03788_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08189__A2 (.I(_03788_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08467__A2 (.I(_03790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08347__A2 (.I(_03790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08267__A2 (.I(_03790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08257__A2 (.I(_03790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08250__A2 (.I(_03790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08244__A2 (.I(_03790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08234__A2 (.I(_03790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08223__B (.I(_03790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08192__A2 (.I(_03790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08512__B2 (.I(_03791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08501__C (.I(_03791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08325__B (.I(_03791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08280__A1 (.I(_03791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08224__A1 (.I(_03791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08192__B (.I(_03791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08194__A2 (.I(_03793_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08404__A2 (.I(_03796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08335__A1 (.I(_03796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08286__A1 (.I(_03796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08217__A1 (.I(_03796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08198__I (.I(_03796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09560__A1 (.I(_03797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08831__S (.I(_03797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08802__A2 (.I(_03797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08514__A1 (.I(_03797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08503__C (.I(_03797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08494__C (.I(_03797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08484__C (.I(_03797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08455__A2 (.I(_03797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08452__A2 (.I(_03797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08442__B (.I(_03797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08379__A1 (.I(_03797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08374__A1 (.I(_03797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08354__C (.I(_03797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08344__B (.I(_03797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08225__C (.I(_03797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08199__I (.I(_03797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09395__A2 (.I(_03798_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08919__A2 (.I(_03798_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08837__A2 (.I(_03798_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08820__A2 (.I(_03798_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08812__B2 (.I(_03798_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08521__A1 (.I(_03798_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08520__A2 (.I(_03798_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08472__A2 (.I(_03798_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08458__A3 (.I(_03798_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08449__A2 (.I(_03798_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08444__B2 (.I(_03798_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08337__A2 (.I(_03798_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08226__A2 (.I(_03798_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08219__A2 (.I(_03798_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08208__A1 (.I(_03798_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08207__A2 (.I(_03798_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08389__C (.I(_03800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08370__B1 (.I(_03800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08327__C (.I(_03800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08273__A1 (.I(_03800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08259__A2 (.I(_03800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08255__C (.I(_03800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08210__A2 (.I(_03800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08202__A2 (.I(_03800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08828__A1 (.I(_03801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08477__B (.I(_03801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08468__C (.I(_03801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08460__B (.I(_03801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08437__C (.I(_03801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08278__A1 (.I(_03801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08251__B1 (.I(_03801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08245__B1 (.I(_03801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08238__B2 (.I(_03801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08205__A1 (.I(_03801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08418__A1 (.I(_03802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08270__A2 (.I(_03802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08246__A2 (.I(_03802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08234__C2 (.I(_03802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08221__A2 (.I(_03802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08204__A2 (.I(_03802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08834__B (.I(_03807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08431__A1 (.I(_03807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08210__A3 (.I(_03807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08835__A2 (.I(_03809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08815__B1 (.I(_03809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08431__A2 (.I(_03809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08256__A3 (.I(_03809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08212__A2 (.I(_03809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08817__A1 (.I(_03810_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08388__A2 (.I(_03810_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08367__A1 (.I(_03810_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08223__C (.I(_03810_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08215__A2 (.I(_03810_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09396__A1 (.I(_03812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08819__A1 (.I(_03812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08403__A1 (.I(_03812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08392__A1 (.I(_03812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08215__B (.I(_03812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08812__A2 (.I(_03816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08520__B1 (.I(_03816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08441__A2 (.I(_03816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08421__A1 (.I(_03816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08414__A1 (.I(_03816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08406__A1 (.I(_03816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08393__C2 (.I(_03816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08377__A1 (.I(_03816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08363__C2 (.I(_03816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08308__A1 (.I(_03816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08287__A1 (.I(_03816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08275__A1 (.I(_03816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08263__A1 (.I(_03816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08229__B1 (.I(_03816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08219__B2 (.I(_03816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08804__A2 (.I(_03818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08479__A2 (.I(_03818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08436__A2 (.I(_03818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08417__C (.I(_03818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08347__B1 (.I(_03818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08250__B1 (.I(_03818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08242__A2 (.I(_03818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08234__B1 (.I(_03818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08223__A1 (.I(_03818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08821__A1 (.I(_03825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08807__A2 (.I(_03825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08481__A2 (.I(_03825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08463__A1 (.I(_03825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08281__A1 (.I(_03825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08238__A1 (.I(_03825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08816__A2 (.I(_03826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08418__A2 (.I(_03826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08402__A3 (.I(_03826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08351__C (.I(_03826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08329__C1 (.I(_03826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08238__A2 (.I(_03826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08479__A1 (.I(_03828_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08434__A2 (.I(_03828_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08398__B1 (.I(_03828_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08389__B1 (.I(_03828_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08327__B1 (.I(_03828_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08324__B1 (.I(_03828_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08283__A2 (.I(_03828_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08266__A2 (.I(_03828_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08260__A2 (.I(_03828_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08234__C1 (.I(_03828_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08434__A1 (.I(_03831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08432__A2 (.I(_03831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08398__B2 (.I(_03831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08370__A1 (.I(_03831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08368__A1 (.I(_03831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08347__A1 (.I(_03831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08325__A1 (.I(_03831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08320__A2 (.I(_03831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08317__A1 (.I(_03831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08312__A1 (.I(_03831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08267__A1 (.I(_03831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08257__B (.I(_03831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08237__B (.I(_03831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08453__B2 (.I(_03834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08240__B (.I(_03834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08518__A1 (.I(_03835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08466__A1 (.I(_03835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08250__C (.I(_03835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08244__B (.I(_03835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08456__B2 (.I(_03840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08247__B (.I(_03840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08834__C (.I(_03851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08826__C (.I(_03851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08493__C (.I(_03851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08489__C (.I(_03851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08481__B (.I(_03851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08476__B (.I(_03851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08465__A1 (.I(_03851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08439__C (.I(_03851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08409__A2 (.I(_03851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08402__A2 (.I(_03851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08391__C (.I(_03851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08353__A1 (.I(_03851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08352__B (.I(_03851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08285__A1 (.I(_03851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08284__C (.I(_03851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08260__B (.I(_03851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08263__B (.I(_03854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08450__B2 (.I(_03855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08339__C (.I(_03855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08264__B (.I(_03855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08275__A2 (.I(_03856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08804__A1 (.I(_03860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08500__A2 (.I(_03860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08389__A2 (.I(_03860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08386__A2 (.I(_03860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08327__A2 (.I(_03860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08272__A2 (.I(_03860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08342__A1 (.I(_03866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08276__B (.I(_03866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08287__A2 (.I(_03867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08284__B2 (.I(_03867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08441__B2 (.I(_03876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08371__A1 (.I(_03876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08362__A1 (.I(_03876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08331__C (.I(_03876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08287__B2 (.I(_03876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08345__B2 (.I(_03877_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08288__B (.I(_03877_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08306__A2 (.I(_03879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08305__A2 (.I(_03879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08304__A2 (.I(_03879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08303__A2 (.I(_03879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08302__A2 (.I(_03879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08301__A2 (.I(_03879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08300__A2 (.I(_03879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08299__A2 (.I(_03879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08298__A2 (.I(_03879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08297__A2 (.I(_03879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08296__A2 (.I(_03879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08295__A2 (.I(_03879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08294__A2 (.I(_03879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08293__A2 (.I(_03879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08292__A2 (.I(_03879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08291__A2 (.I(_03879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08467__A1 (.I(_03890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08352__A1 (.I(_03890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08329__A2 (.I(_03890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08324__B2 (.I(_03890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08314__A1 (.I(_03890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08476__C (.I(_03896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08465__A2 (.I(_03896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08391__A2 (.I(_03896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08352__A2 (.I(_03896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08316__A2 (.I(_03896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08817__B (.I(_03897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08805__A2 (.I(_03897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08501__A2 (.I(_03897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08491__A2 (.I(_03897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08411__A1 (.I(_03897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08325__A2 (.I(_03897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08323__A1 (.I(_03897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08521__A2 (.I(_03906_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08420__B (.I(_03906_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08411__B (.I(_03906_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08399__B (.I(_03906_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08326__B (.I(_03906_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08384__A1 (.I(_03913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08333__B (.I(_03913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08344__A2 (.I(_03914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08340__A2 (.I(_03914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08335__A2 (.I(_03914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08363__A2 (.I(_03916_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08357__A1 (.I(_03916_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08356__A2 (.I(_03916_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08345__A2 (.I(_03916_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08341__A2 (.I(_03916_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08339__A1 (.I(_03916_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08338__A2 (.I(_03916_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08354__A2 (.I(_03923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08351__A2 (.I(_03923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08353__A2 (.I(_03926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08357__A2 (.I(_03931_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08363__C1 (.I(_03935_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08360__B2 (.I(_03935_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08482__C (.I(_03940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08370__B2 (.I(_03940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08404__A3 (.I(_03947_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08373__A2 (.I(_03947_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08393__C1 (.I(_03963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08391__B1 (.I(_03963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08394__A1 (.I(_03965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08823__A1 (.I(_03973_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08815__A1 (.I(_03973_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08493__A1 (.I(_03973_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08460__A1 (.I(_03973_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08402__A1 (.I(_03973_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08406__B (.I(_03975_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08414__B (.I(_03983_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08421__A2 (.I(_03985_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08420__A1 (.I(_03987_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08518__A2 (.I(_03988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08507__A2 (.I(_03988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08477__A2 (.I(_03988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08468__A2 (.I(_03988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08466__A2 (.I(_03988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08460__A2 (.I(_03988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08437__A2 (.I(_03988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08419__B (.I(_03988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08920__A1 (.I(_03991_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08428__A1 (.I(_03991_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08470__A1 (.I(_03999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08468__A1 (.I(_03999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08437__A1 (.I(_03999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08435__A1 (.I(_03999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08433__A1 (.I(_03999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08441__B1 (.I(_04009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08803__B2 (.I(_04010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08444__A1 (.I(_04010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08517__A1 (.I(_04016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08516__A2 (.I(_04016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08506__A1 (.I(_04016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08505__A2 (.I(_04016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08497__A1 (.I(_04016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08496__A2 (.I(_04016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08487__A1 (.I(_04016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08486__A2 (.I(_04016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08473__A2 (.I(_04016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08472__B (.I(_04016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08457__A2 (.I(_04016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08456__A2 (.I(_04016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08453__A2 (.I(_04016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08452__B (.I(_04016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08450__A2 (.I(_04016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08449__B (.I(_04016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08818__B2 (.I(_04024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08492__A1 (.I(_04024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08464__A1 (.I(_04024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08473__B1 (.I(_04035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08480__A2 (.I(_04041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08503__A2 (.I(_04059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08511__A2 (.I(_04070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08517__A3 (.I(_04075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08520__B2 (.I(_04078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08543__A2 (.I(_04084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08542__A2 (.I(_04084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08541__A2 (.I(_04084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08540__A2 (.I(_04084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08539__A2 (.I(_04084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08538__A2 (.I(_04084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08537__A2 (.I(_04084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08536__A2 (.I(_04084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08535__A2 (.I(_04084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08534__A2 (.I(_04084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08533__A2 (.I(_04084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08532__A2 (.I(_04084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08531__A2 (.I(_04084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08530__A2 (.I(_04084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08529__A2 (.I(_04084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08528__A2 (.I(_04084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08561__A2 (.I(_04094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08560__A2 (.I(_04094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08559__A2 (.I(_04094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08558__A2 (.I(_04094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08557__A2 (.I(_04094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08556__A2 (.I(_04094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08555__A2 (.I(_04094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08554__A2 (.I(_04094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08553__A2 (.I(_04094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08552__A2 (.I(_04094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08551__A2 (.I(_04094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08550__A2 (.I(_04094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08549__A2 (.I(_04094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08548__A2 (.I(_04094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08547__A2 (.I(_04094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08546__A2 (.I(_04094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08617__S (.I(_04115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08615__S (.I(_04115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08613__S (.I(_04115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08611__S (.I(_04115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08609__S (.I(_04115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08607__S (.I(_04115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08605__S (.I(_04115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08603__S (.I(_04115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08601__S (.I(_04115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08599__S (.I(_04115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08597__S (.I(_04115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08595__S (.I(_04115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08593__S (.I(_04115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08591__S (.I(_04115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08589__S (.I(_04115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08587__S (.I(_04115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08633__A1 (.I(_04137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08627__B1 (.I(_04137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08653__A2 (.I(_04145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08652__A2 (.I(_04145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08651__A2 (.I(_04145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08650__A2 (.I(_04145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08649__A2 (.I(_04145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08648__A2 (.I(_04145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08647__A2 (.I(_04145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08646__A2 (.I(_04145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08645__A2 (.I(_04145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08644__A2 (.I(_04145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08643__A2 (.I(_04145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08642__A2 (.I(_04145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08641__A2 (.I(_04145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08640__A2 (.I(_04145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08639__A2 (.I(_04145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08638__A2 (.I(_04145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09562__A1 (.I(_04155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08686__A2 (.I(_04155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08684__A2 (.I(_04155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08682__A2 (.I(_04155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08680__A2 (.I(_04155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08678__A2 (.I(_04155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08676__A2 (.I(_04155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08674__A2 (.I(_04155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08672__A2 (.I(_04155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08670__A2 (.I(_04155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08668__A2 (.I(_04155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08666__A2 (.I(_04155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08664__A2 (.I(_04155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08662__A2 (.I(_04155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08660__A2 (.I(_04155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08658__A2 (.I(_04155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08689__B1 (.I(_04157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08686__B1 (.I(_04157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08684__B1 (.I(_04157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08682__B1 (.I(_04157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08680__B1 (.I(_04157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08678__B1 (.I(_04157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08676__B1 (.I(_04157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08674__B1 (.I(_04157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08672__B1 (.I(_04157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08670__B1 (.I(_04157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08668__B1 (.I(_04157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08666__B1 (.I(_04157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08664__B1 (.I(_04157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08662__B1 (.I(_04157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08660__B1 (.I(_04157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08658__B1 (.I(_04157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08720__A2 (.I(_04173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08718__A2 (.I(_04173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08716__A2 (.I(_04173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08714__A2 (.I(_04173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08712__A2 (.I(_04173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08710__A2 (.I(_04173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08708__A2 (.I(_04173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08706__A2 (.I(_04173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08704__A2 (.I(_04173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08702__A2 (.I(_04173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08700__A2 (.I(_04173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08698__A2 (.I(_04173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08696__A2 (.I(_04173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08694__A2 (.I(_04173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08692__A2 (.I(_04173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08689__A2 (.I(_04173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08727__B1 (.I(_04175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08720__B1 (.I(_04175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08718__B1 (.I(_04175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08716__B1 (.I(_04175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08714__B1 (.I(_04175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08712__B1 (.I(_04175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08710__B1 (.I(_04175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08708__B1 (.I(_04175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08706__B1 (.I(_04175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08704__B1 (.I(_04175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08702__B1 (.I(_04175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08700__B1 (.I(_04175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08698__B1 (.I(_04175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08696__B1 (.I(_04175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08694__B1 (.I(_04175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08692__B1 (.I(_04175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09392__A1 (.I(_04191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09390__A1 (.I(_04191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08723__A1 (.I(_04191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08727__B2 (.I(_04195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09506__A2 (.I(_04197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09488__A2 (.I(_04197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09306__A2 (.I(_04197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09270__A2 (.I(_04197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09155__A2 (.I(_04197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09119__A2 (.I(_04197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09101__A2 (.I(_04197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09083__A2 (.I(_04197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09047__A2 (.I(_04197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09029__A2 (.I(_04197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09011__A2 (.I(_04197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08993__A2 (.I(_04197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08975__A2 (.I(_04197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08901__A2 (.I(_04197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08839__A2 (.I(_04197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08730__A2 (.I(_04197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08747__A2 (.I(_04199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08746__A2 (.I(_04199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08745__A2 (.I(_04199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08744__A2 (.I(_04199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08743__A2 (.I(_04199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08742__A2 (.I(_04199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08741__A2 (.I(_04199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08740__A2 (.I(_04199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08739__A2 (.I(_04199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08738__A2 (.I(_04199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08737__A2 (.I(_04199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08736__A2 (.I(_04199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08735__A2 (.I(_04199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08734__A2 (.I(_04199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08733__A2 (.I(_04199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08732__A2 (.I(_04199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08763__S (.I(_04208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08761__S (.I(_04208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08759__S (.I(_04208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08757__S (.I(_04208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08755__S (.I(_04208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08753__S (.I(_04208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08751__S (.I(_04208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08749__S (.I(_04208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08780__S (.I(_04217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08778__S (.I(_04217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08776__S (.I(_04217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08774__S (.I(_04217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08772__S (.I(_04217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08770__S (.I(_04217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08768__S (.I(_04217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08766__S (.I(_04217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08799__A2 (.I(_04227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08798__A2 (.I(_04227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08797__A2 (.I(_04227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08796__A2 (.I(_04227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08795__A2 (.I(_04227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08794__A2 (.I(_04227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08793__A2 (.I(_04227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08792__A2 (.I(_04227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08791__A2 (.I(_04227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08790__A2 (.I(_04227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08789__A2 (.I(_04227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08788__A2 (.I(_04227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08787__A2 (.I(_04227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08786__A2 (.I(_04227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08785__A2 (.I(_04227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08784__A2 (.I(_04227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08810__A2 (.I(_04242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08856__A2 (.I(_04271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08855__A2 (.I(_04271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08854__A2 (.I(_04271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08853__A2 (.I(_04271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08852__A2 (.I(_04271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08851__A2 (.I(_04271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08850__A2 (.I(_04271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08849__A2 (.I(_04271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08848__A2 (.I(_04271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08847__A2 (.I(_04271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08846__A2 (.I(_04271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08845__A2 (.I(_04271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08844__A2 (.I(_04271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08843__A2 (.I(_04271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08842__A2 (.I(_04271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08841__A2 (.I(_04271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09176__A1 (.I(_04280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09158__A1 (.I(_04280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09140__A1 (.I(_04280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09122__A1 (.I(_04280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09104__A1 (.I(_04280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09086__A1 (.I(_04280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09068__A1 (.I(_04280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09050__A1 (.I(_04280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09032__A1 (.I(_04280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09014__A1 (.I(_04280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08996__A1 (.I(_04280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08978__A1 (.I(_04280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08927__A1 (.I(_04280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08904__A1 (.I(_04280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08886__A1 (.I(_04280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08861__A1 (.I(_04280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08882__A2 (.I(_04282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08881__A2 (.I(_04282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08879__A2 (.I(_04282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08878__A2 (.I(_04282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08876__A2 (.I(_04282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08875__A2 (.I(_04282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08873__A2 (.I(_04282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08872__A2 (.I(_04282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08870__A2 (.I(_04282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08869__A2 (.I(_04282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08867__A2 (.I(_04282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08866__A2 (.I(_04282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08864__A2 (.I(_04282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08863__A2 (.I(_04282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08861__A2 (.I(_04282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08860__A2 (.I(_04282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09178__A1 (.I(_04284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09160__A1 (.I(_04284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09142__A1 (.I(_04284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09124__A1 (.I(_04284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09106__A1 (.I(_04284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09088__A1 (.I(_04284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09070__A1 (.I(_04284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09052__A1 (.I(_04284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09034__A1 (.I(_04284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09016__A1 (.I(_04284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08998__A1 (.I(_04284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08980__A1 (.I(_04284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08929__A1 (.I(_04284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08906__A1 (.I(_04284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08888__A1 (.I(_04284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08864__A1 (.I(_04284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09180__A1 (.I(_04286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09162__A1 (.I(_04286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09144__A1 (.I(_04286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09126__A1 (.I(_04286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09108__A1 (.I(_04286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09090__A1 (.I(_04286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09072__A1 (.I(_04286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09054__A1 (.I(_04286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09036__A1 (.I(_04286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09018__A1 (.I(_04286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09000__A1 (.I(_04286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08982__A1 (.I(_04286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08931__A1 (.I(_04286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08908__A1 (.I(_04286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08890__A1 (.I(_04286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08867__A1 (.I(_04286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09182__A1 (.I(_04288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09164__A1 (.I(_04288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09146__A1 (.I(_04288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09128__A1 (.I(_04288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09110__A1 (.I(_04288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09092__A1 (.I(_04288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09074__A1 (.I(_04288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09056__A1 (.I(_04288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09038__A1 (.I(_04288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09020__A1 (.I(_04288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09002__A1 (.I(_04288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08984__A1 (.I(_04288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08933__A1 (.I(_04288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08910__A1 (.I(_04288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08892__A1 (.I(_04288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08870__A1 (.I(_04288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09184__A1 (.I(_04290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09166__A1 (.I(_04290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09148__A1 (.I(_04290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09130__A1 (.I(_04290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09112__A1 (.I(_04290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09094__A1 (.I(_04290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09076__A1 (.I(_04290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09058__A1 (.I(_04290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09040__A1 (.I(_04290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09022__A1 (.I(_04290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09004__A1 (.I(_04290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08986__A1 (.I(_04290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08935__A1 (.I(_04290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08912__A1 (.I(_04290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08894__A1 (.I(_04290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08873__A1 (.I(_04290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09186__A1 (.I(_04292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09168__A1 (.I(_04292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09150__A1 (.I(_04292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09132__A1 (.I(_04292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09114__A1 (.I(_04292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09096__A1 (.I(_04292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09078__A1 (.I(_04292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09060__A1 (.I(_04292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09042__A1 (.I(_04292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09024__A1 (.I(_04292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09006__A1 (.I(_04292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08988__A1 (.I(_04292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08937__A1 (.I(_04292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08914__A1 (.I(_04292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08896__A1 (.I(_04292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08876__A1 (.I(_04292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09188__A1 (.I(_04294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09170__A1 (.I(_04294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09152__A1 (.I(_04294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09134__A1 (.I(_04294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09116__A1 (.I(_04294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09098__A1 (.I(_04294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09080__A1 (.I(_04294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09062__A1 (.I(_04294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09044__A1 (.I(_04294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09026__A1 (.I(_04294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09008__A1 (.I(_04294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08990__A1 (.I(_04294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08939__A1 (.I(_04294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08916__A1 (.I(_04294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08898__A1 (.I(_04294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08879__A1 (.I(_04294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09190__A1 (.I(_04296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09172__A1 (.I(_04296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09154__A1 (.I(_04296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09136__A1 (.I(_04296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09118__A1 (.I(_04296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09100__A1 (.I(_04296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09082__A1 (.I(_04296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09064__A1 (.I(_04296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09046__A1 (.I(_04296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09028__A1 (.I(_04296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09010__A1 (.I(_04296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08992__A1 (.I(_04296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08941__A1 (.I(_04296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08918__A1 (.I(_04296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08900__A1 (.I(_04296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08882__A1 (.I(_04296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08900__A2 (.I(_04299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08899__A2 (.I(_04299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08898__A2 (.I(_04299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08897__A2 (.I(_04299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08896__A2 (.I(_04299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08895__A2 (.I(_04299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08894__A2 (.I(_04299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08893__A2 (.I(_04299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08892__A2 (.I(_04299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08891__A2 (.I(_04299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08890__A2 (.I(_04299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08889__A2 (.I(_04299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08888__A2 (.I(_04299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08887__A2 (.I(_04299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08886__A2 (.I(_04299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08885__A2 (.I(_04299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08918__A2 (.I(_04309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08917__A2 (.I(_04309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08916__A2 (.I(_04309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08915__A2 (.I(_04309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08914__A2 (.I(_04309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08913__A2 (.I(_04309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08912__A2 (.I(_04309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08911__A2 (.I(_04309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08910__A2 (.I(_04309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08909__A2 (.I(_04309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08908__A2 (.I(_04309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08907__A2 (.I(_04309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08906__A2 (.I(_04309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08905__A2 (.I(_04309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08904__A2 (.I(_04309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08903__A2 (.I(_04309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08941__A2 (.I(_04322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08940__A2 (.I(_04322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08939__A2 (.I(_04322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08938__A2 (.I(_04322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08937__A2 (.I(_04322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08936__A2 (.I(_04322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08935__A2 (.I(_04322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08934__A2 (.I(_04322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08933__A2 (.I(_04322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08932__A2 (.I(_04322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08931__A2 (.I(_04322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08930__A2 (.I(_04322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08929__A2 (.I(_04322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08928__A2 (.I(_04322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08927__A2 (.I(_04322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08926__A2 (.I(_04322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08973__S (.I(_04331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08971__S (.I(_04331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08969__S (.I(_04331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08967__S (.I(_04331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08965__S (.I(_04331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08963__S (.I(_04331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08961__S (.I(_04331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08959__S (.I(_04331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08957__S (.I(_04331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08955__S (.I(_04331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08953__S (.I(_04331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08951__S (.I(_04331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08949__S (.I(_04331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08947__S (.I(_04331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08945__S (.I(_04331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08943__S (.I(_04331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08992__A2 (.I(_04349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08991__A2 (.I(_04349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08990__A2 (.I(_04349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08989__A2 (.I(_04349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08988__A2 (.I(_04349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08987__A2 (.I(_04349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08986__A2 (.I(_04349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08985__A2 (.I(_04349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08984__A2 (.I(_04349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08983__A2 (.I(_04349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08982__A2 (.I(_04349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08981__A2 (.I(_04349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08980__A2 (.I(_04349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08979__A2 (.I(_04349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08978__A2 (.I(_04349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08977__A2 (.I(_04349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09010__A2 (.I(_04359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09009__A2 (.I(_04359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09008__A2 (.I(_04359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09007__A2 (.I(_04359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09006__A2 (.I(_04359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09005__A2 (.I(_04359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09004__A2 (.I(_04359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09003__A2 (.I(_04359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09002__A2 (.I(_04359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09001__A2 (.I(_04359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09000__A2 (.I(_04359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08999__A2 (.I(_04359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08998__A2 (.I(_04359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08997__A2 (.I(_04359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08996__A2 (.I(_04359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08995__A2 (.I(_04359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09028__A2 (.I(_04369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09027__A2 (.I(_04369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09026__A2 (.I(_04369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09025__A2 (.I(_04369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09024__A2 (.I(_04369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09023__A2 (.I(_04369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09022__A2 (.I(_04369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09021__A2 (.I(_04369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09020__A2 (.I(_04369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09019__A2 (.I(_04369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09018__A2 (.I(_04369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09017__A2 (.I(_04369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09016__A2 (.I(_04369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09015__A2 (.I(_04369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09014__A2 (.I(_04369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09013__A2 (.I(_04369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09046__A2 (.I(_04379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09045__A2 (.I(_04379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09044__A2 (.I(_04379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09043__A2 (.I(_04379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09042__A2 (.I(_04379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09041__A2 (.I(_04379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09040__A2 (.I(_04379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09039__A2 (.I(_04379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09038__A2 (.I(_04379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09037__A2 (.I(_04379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09036__A2 (.I(_04379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09035__A2 (.I(_04379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09034__A2 (.I(_04379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09033__A2 (.I(_04379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09032__A2 (.I(_04379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09031__A2 (.I(_04379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09064__A2 (.I(_04389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09063__A2 (.I(_04389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09062__A2 (.I(_04389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09061__A2 (.I(_04389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09060__A2 (.I(_04389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09059__A2 (.I(_04389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09058__A2 (.I(_04389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09057__A2 (.I(_04389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09056__A2 (.I(_04389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09055__A2 (.I(_04389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09054__A2 (.I(_04389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09053__A2 (.I(_04389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09052__A2 (.I(_04389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09051__A2 (.I(_04389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09050__A2 (.I(_04389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09049__A2 (.I(_04389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09082__A2 (.I(_04399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09081__A2 (.I(_04399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09080__A2 (.I(_04399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09079__A2 (.I(_04399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09078__A2 (.I(_04399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09077__A2 (.I(_04399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09076__A2 (.I(_04399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09075__A2 (.I(_04399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09074__A2 (.I(_04399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09073__A2 (.I(_04399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09072__A2 (.I(_04399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09071__A2 (.I(_04399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09070__A2 (.I(_04399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09069__A2 (.I(_04399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09068__A2 (.I(_04399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09067__A2 (.I(_04399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09100__A2 (.I(_04409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09099__A2 (.I(_04409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09098__A2 (.I(_04409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09097__A2 (.I(_04409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09096__A2 (.I(_04409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09095__A2 (.I(_04409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09094__A2 (.I(_04409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09093__A2 (.I(_04409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09092__A2 (.I(_04409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09091__A2 (.I(_04409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09090__A2 (.I(_04409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09089__A2 (.I(_04409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09088__A2 (.I(_04409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09087__A2 (.I(_04409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09086__A2 (.I(_04409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09085__A2 (.I(_04409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09118__A2 (.I(_04419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09117__A2 (.I(_04419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09116__A2 (.I(_04419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09115__A2 (.I(_04419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09114__A2 (.I(_04419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09113__A2 (.I(_04419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09112__A2 (.I(_04419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09111__A2 (.I(_04419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09110__A2 (.I(_04419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09109__A2 (.I(_04419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09108__A2 (.I(_04419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09107__A2 (.I(_04419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09106__A2 (.I(_04419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09105__A2 (.I(_04419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09104__A2 (.I(_04419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09103__A2 (.I(_04419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09136__A2 (.I(_04429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09135__A2 (.I(_04429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09134__A2 (.I(_04429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09133__A2 (.I(_04429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09132__A2 (.I(_04429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09131__A2 (.I(_04429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09130__A2 (.I(_04429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09129__A2 (.I(_04429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09128__A2 (.I(_04429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09127__A2 (.I(_04429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09126__A2 (.I(_04429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09125__A2 (.I(_04429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09124__A2 (.I(_04429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09123__A2 (.I(_04429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09122__A2 (.I(_04429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09121__A2 (.I(_04429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09154__A2 (.I(_04439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09153__A2 (.I(_04439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09152__A2 (.I(_04439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09151__A2 (.I(_04439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09150__A2 (.I(_04439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09149__A2 (.I(_04439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09148__A2 (.I(_04439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09147__A2 (.I(_04439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09146__A2 (.I(_04439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09145__A2 (.I(_04439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09144__A2 (.I(_04439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09143__A2 (.I(_04439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09142__A2 (.I(_04439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09141__A2 (.I(_04439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09140__A2 (.I(_04439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09139__A2 (.I(_04439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09172__A2 (.I(_04449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09171__A2 (.I(_04449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09170__A2 (.I(_04449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09169__A2 (.I(_04449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09168__A2 (.I(_04449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09167__A2 (.I(_04449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09166__A2 (.I(_04449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09165__A2 (.I(_04449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09164__A2 (.I(_04449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09163__A2 (.I(_04449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09162__A2 (.I(_04449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09161__A2 (.I(_04449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09160__A2 (.I(_04449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09159__A2 (.I(_04449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09158__A2 (.I(_04449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09157__A2 (.I(_04449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09190__A2 (.I(_04459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09189__A2 (.I(_04459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09188__A2 (.I(_04459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09187__A2 (.I(_04459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09186__A2 (.I(_04459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09185__A2 (.I(_04459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09184__A2 (.I(_04459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09183__A2 (.I(_04459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09182__A2 (.I(_04459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09181__A2 (.I(_04459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09180__A2 (.I(_04459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09179__A2 (.I(_04459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09178__A2 (.I(_04459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09177__A2 (.I(_04459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09176__A2 (.I(_04459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09175__A2 (.I(_04459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09545__A1 (.I(_04468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09527__A1 (.I(_04468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09509__A1 (.I(_04468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09491__A1 (.I(_04468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09456__A1 (.I(_04468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09438__A1 (.I(_04468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09420__A1 (.I(_04468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09402__A1 (.I(_04468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09345__A1 (.I(_04468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09327__A1 (.I(_04468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09309__A1 (.I(_04468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09291__A1 (.I(_04468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09273__A1 (.I(_04468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09255__A1 (.I(_04468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09220__A1 (.I(_04468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09195__A1 (.I(_04468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09216__A2 (.I(_04470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09215__A2 (.I(_04470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09213__A2 (.I(_04470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09212__A2 (.I(_04470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09210__A2 (.I(_04470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09209__A2 (.I(_04470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09207__A2 (.I(_04470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09206__A2 (.I(_04470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09204__A2 (.I(_04470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09203__A2 (.I(_04470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09201__A2 (.I(_04470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09200__A2 (.I(_04470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09198__A2 (.I(_04470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09197__A2 (.I(_04470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09195__A2 (.I(_04470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09194__A2 (.I(_04470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09547__A1 (.I(_04472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09529__A1 (.I(_04472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09511__A1 (.I(_04472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09493__A1 (.I(_04472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09458__A1 (.I(_04472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09440__A1 (.I(_04472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09422__A1 (.I(_04472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09404__A1 (.I(_04472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09347__A1 (.I(_04472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09329__A1 (.I(_04472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09311__A1 (.I(_04472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09293__A1 (.I(_04472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09275__A1 (.I(_04472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09257__A1 (.I(_04472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09222__A1 (.I(_04472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09198__A1 (.I(_04472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09549__A1 (.I(_04474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09531__A1 (.I(_04474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09513__A1 (.I(_04474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09495__A1 (.I(_04474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09460__A1 (.I(_04474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09442__A1 (.I(_04474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09424__A1 (.I(_04474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09406__A1 (.I(_04474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09349__A1 (.I(_04474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09331__A1 (.I(_04474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09313__A1 (.I(_04474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09295__A1 (.I(_04474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09277__A1 (.I(_04474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09259__A1 (.I(_04474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09224__A1 (.I(_04474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09201__A1 (.I(_04474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09551__A1 (.I(_04476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09533__A1 (.I(_04476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09515__A1 (.I(_04476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09497__A1 (.I(_04476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09462__A1 (.I(_04476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09444__A1 (.I(_04476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09426__A1 (.I(_04476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09408__A1 (.I(_04476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09351__A1 (.I(_04476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09333__A1 (.I(_04476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09315__A1 (.I(_04476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09297__A1 (.I(_04476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09279__A1 (.I(_04476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09261__A1 (.I(_04476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09226__A1 (.I(_04476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09204__A1 (.I(_04476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09553__A1 (.I(_04478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09535__A1 (.I(_04478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09517__A1 (.I(_04478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09499__A1 (.I(_04478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09464__A1 (.I(_04478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09446__A1 (.I(_04478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09428__A1 (.I(_04478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09410__A1 (.I(_04478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09353__A1 (.I(_04478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09335__A1 (.I(_04478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09317__A1 (.I(_04478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09299__A1 (.I(_04478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09281__A1 (.I(_04478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09263__A1 (.I(_04478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09228__A1 (.I(_04478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09207__A1 (.I(_04478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09555__A1 (.I(_04480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09537__A1 (.I(_04480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09519__A1 (.I(_04480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09501__A1 (.I(_04480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09466__A1 (.I(_04480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09448__A1 (.I(_04480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09430__A1 (.I(_04480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09412__A1 (.I(_04480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09355__A1 (.I(_04480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09337__A1 (.I(_04480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09319__A1 (.I(_04480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09301__A1 (.I(_04480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09283__A1 (.I(_04480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09265__A1 (.I(_04480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09230__A1 (.I(_04480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09210__A1 (.I(_04480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09557__A1 (.I(_04482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09539__A1 (.I(_04482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09521__A1 (.I(_04482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09503__A1 (.I(_04482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09468__A1 (.I(_04482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09450__A1 (.I(_04482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09432__A1 (.I(_04482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09414__A1 (.I(_04482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09357__A1 (.I(_04482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09339__A1 (.I(_04482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09321__A1 (.I(_04482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09303__A1 (.I(_04482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09285__A1 (.I(_04482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09267__A1 (.I(_04482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09232__A1 (.I(_04482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09213__A1 (.I(_04482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09559__A1 (.I(_04484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09541__A1 (.I(_04484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09523__A1 (.I(_04484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09505__A1 (.I(_04484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09470__A1 (.I(_04484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09452__A1 (.I(_04484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09434__A1 (.I(_04484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09416__A1 (.I(_04484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09359__A1 (.I(_04484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09341__A1 (.I(_04484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09323__A1 (.I(_04484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09305__A1 (.I(_04484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09287__A1 (.I(_04484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09269__A1 (.I(_04484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09234__A1 (.I(_04484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09216__A1 (.I(_04484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09234__A2 (.I(_04487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09233__A2 (.I(_04487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09232__A2 (.I(_04487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09231__A2 (.I(_04487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09230__A2 (.I(_04487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09229__A2 (.I(_04487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09228__A2 (.I(_04487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09227__A2 (.I(_04487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09226__A2 (.I(_04487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09225__A2 (.I(_04487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09224__A2 (.I(_04487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09223__A2 (.I(_04487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09222__A2 (.I(_04487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09221__A2 (.I(_04487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09220__A2 (.I(_04487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09219__A2 (.I(_04487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09250__S (.I(_04496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09248__S (.I(_04496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09246__S (.I(_04496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09244__S (.I(_04496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09242__S (.I(_04496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09240__S (.I(_04496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09238__S (.I(_04496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09236__S (.I(_04496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09269__A2 (.I(_04506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09268__A2 (.I(_04506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09267__A2 (.I(_04506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09266__A2 (.I(_04506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09265__A2 (.I(_04506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09264__A2 (.I(_04506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09263__A2 (.I(_04506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09262__A2 (.I(_04506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09261__A2 (.I(_04506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09260__A2 (.I(_04506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09259__A2 (.I(_04506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09258__A2 (.I(_04506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09257__A2 (.I(_04506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09256__A2 (.I(_04506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09255__A2 (.I(_04506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09254__A2 (.I(_04506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09287__A2 (.I(_04516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09286__A2 (.I(_04516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09285__A2 (.I(_04516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09284__A2 (.I(_04516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09283__A2 (.I(_04516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09282__A2 (.I(_04516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09281__A2 (.I(_04516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09280__A2 (.I(_04516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09279__A2 (.I(_04516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09278__A2 (.I(_04516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09277__A2 (.I(_04516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09276__A2 (.I(_04516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09275__A2 (.I(_04516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09274__A2 (.I(_04516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09273__A2 (.I(_04516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09272__A2 (.I(_04516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09305__A2 (.I(_04526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09304__A2 (.I(_04526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09303__A2 (.I(_04526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09302__A2 (.I(_04526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09301__A2 (.I(_04526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09300__A2 (.I(_04526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09299__A2 (.I(_04526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09298__A2 (.I(_04526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09297__A2 (.I(_04526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09296__A2 (.I(_04526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09295__A2 (.I(_04526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09294__A2 (.I(_04526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09293__A2 (.I(_04526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09292__A2 (.I(_04526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09291__A2 (.I(_04526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09290__A2 (.I(_04526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09323__A2 (.I(_04536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09322__A2 (.I(_04536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09321__A2 (.I(_04536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09320__A2 (.I(_04536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09319__A2 (.I(_04536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09318__A2 (.I(_04536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09317__A2 (.I(_04536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09316__A2 (.I(_04536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09315__A2 (.I(_04536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09314__A2 (.I(_04536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09313__A2 (.I(_04536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09312__A2 (.I(_04536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09311__A2 (.I(_04536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09310__A2 (.I(_04536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09309__A2 (.I(_04536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09308__A2 (.I(_04536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09341__A2 (.I(_04546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09340__A2 (.I(_04546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09339__A2 (.I(_04546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09338__A2 (.I(_04546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09337__A2 (.I(_04546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09336__A2 (.I(_04546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09335__A2 (.I(_04546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09334__A2 (.I(_04546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09333__A2 (.I(_04546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09332__A2 (.I(_04546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09331__A2 (.I(_04546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09330__A2 (.I(_04546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09329__A2 (.I(_04546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09328__A2 (.I(_04546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09327__A2 (.I(_04546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09326__A2 (.I(_04546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09359__A2 (.I(_04556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09358__A2 (.I(_04556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09357__A2 (.I(_04556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09356__A2 (.I(_04556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09355__A2 (.I(_04556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09354__A2 (.I(_04556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09353__A2 (.I(_04556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09352__A2 (.I(_04556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09351__A2 (.I(_04556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09350__A2 (.I(_04556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09349__A2 (.I(_04556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09348__A2 (.I(_04556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09347__A2 (.I(_04556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09346__A2 (.I(_04556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09345__A2 (.I(_04556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09344__A2 (.I(_04556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09378__A2 (.I(_04568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09377__B (.I(_04568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09375__A1 (.I(_04568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09374__A2 (.I(_04568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09371__S (.I(_04568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09368__A2 (.I(_04568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09367__A1 (.I(_04568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09416__A2 (.I(_04595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09415__A2 (.I(_04595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09414__A2 (.I(_04595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09413__A2 (.I(_04595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09412__A2 (.I(_04595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09411__A2 (.I(_04595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09410__A2 (.I(_04595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09409__A2 (.I(_04595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09408__A2 (.I(_04595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09407__A2 (.I(_04595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09406__A2 (.I(_04595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09405__A2 (.I(_04595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09404__A2 (.I(_04595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09403__A2 (.I(_04595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09402__A2 (.I(_04595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09401__A2 (.I(_04595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09434__A2 (.I(_04605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09433__A2 (.I(_04605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09432__A2 (.I(_04605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09431__A2 (.I(_04605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09430__A2 (.I(_04605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09429__A2 (.I(_04605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09428__A2 (.I(_04605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09427__A2 (.I(_04605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09426__A2 (.I(_04605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09425__A2 (.I(_04605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09424__A2 (.I(_04605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09423__A2 (.I(_04605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09422__A2 (.I(_04605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09421__A2 (.I(_04605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09420__A2 (.I(_04605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09419__A2 (.I(_04605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09452__A2 (.I(_04615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09451__A2 (.I(_04615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09450__A2 (.I(_04615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09449__A2 (.I(_04615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09448__A2 (.I(_04615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09447__A2 (.I(_04615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09446__A2 (.I(_04615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09445__A2 (.I(_04615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09444__A2 (.I(_04615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09443__A2 (.I(_04615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09442__A2 (.I(_04615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09441__A2 (.I(_04615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09440__A2 (.I(_04615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09439__A2 (.I(_04615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09438__A2 (.I(_04615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09437__A2 (.I(_04615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09470__A2 (.I(_04625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09469__A2 (.I(_04625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09468__A2 (.I(_04625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09467__A2 (.I(_04625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09466__A2 (.I(_04625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09465__A2 (.I(_04625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09464__A2 (.I(_04625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09463__A2 (.I(_04625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09462__A2 (.I(_04625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09461__A2 (.I(_04625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09460__A2 (.I(_04625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09459__A2 (.I(_04625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09458__A2 (.I(_04625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09457__A2 (.I(_04625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09456__A2 (.I(_04625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09455__A2 (.I(_04625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09486__S (.I(_04634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09484__S (.I(_04634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09482__S (.I(_04634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09480__S (.I(_04634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09478__S (.I(_04634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09476__S (.I(_04634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09474__S (.I(_04634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09472__S (.I(_04634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09505__A2 (.I(_04644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09504__A2 (.I(_04644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09503__A2 (.I(_04644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09502__A2 (.I(_04644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09501__A2 (.I(_04644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09500__A2 (.I(_04644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09499__A2 (.I(_04644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09498__A2 (.I(_04644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09497__A2 (.I(_04644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09496__A2 (.I(_04644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09495__A2 (.I(_04644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09494__A2 (.I(_04644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09493__A2 (.I(_04644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09492__A2 (.I(_04644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09491__A2 (.I(_04644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09490__A2 (.I(_04644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09523__A2 (.I(_04654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09522__A2 (.I(_04654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09521__A2 (.I(_04654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09520__A2 (.I(_04654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09519__A2 (.I(_04654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09518__A2 (.I(_04654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09517__A2 (.I(_04654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09516__A2 (.I(_04654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09515__A2 (.I(_04654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09514__A2 (.I(_04654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09513__A2 (.I(_04654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09512__A2 (.I(_04654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09511__A2 (.I(_04654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09510__A2 (.I(_04654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09509__A2 (.I(_04654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09508__A2 (.I(_04654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09541__A2 (.I(_04664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09540__A2 (.I(_04664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09539__A2 (.I(_04664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09538__A2 (.I(_04664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09537__A2 (.I(_04664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09536__A2 (.I(_04664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09535__A2 (.I(_04664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09534__A2 (.I(_04664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09533__A2 (.I(_04664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09532__A2 (.I(_04664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09531__A2 (.I(_04664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09530__A2 (.I(_04664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09529__A2 (.I(_04664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09528__A2 (.I(_04664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09527__A2 (.I(_04664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09526__A2 (.I(_04664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09559__A2 (.I(_04674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09558__A2 (.I(_04674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09557__A2 (.I(_04674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09556__A2 (.I(_04674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09555__A2 (.I(_04674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09554__A2 (.I(_04674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09553__A2 (.I(_04674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09552__A2 (.I(_04674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09551__A2 (.I(_04674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09550__A2 (.I(_04674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09549__A2 (.I(_04674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09548__A2 (.I(_04674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09547__A2 (.I(_04674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09546__A2 (.I(_04674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09545__A2 (.I(_04674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09544__A2 (.I(_04674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09562__A2 (.I(_04683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09561__A2 (.I(_04683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.input_buf_clk_I  (.I(io_in[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04904__I (.I(io_in[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[0]_D  (.I(io_in[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[25]_SE  (.I(io_in[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[24]_SE  (.I(io_in[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[23]_SE  (.I(io_in[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[22]_SE  (.I(io_in[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[21]_SE  (.I(io_in[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[20]_SE  (.I(io_in[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[19]_SE  (.I(io_in[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[18]_SE  (.I(io_in[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[17]_SE  (.I(io_in[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[16]_SE  (.I(io_in[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[15]_SE  (.I(io_in[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[14]_SE  (.I(io_in[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[26]_SE  (.I(io_in[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[32]_SE  (.I(io_in[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[31]_SE  (.I(io_in[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[27]_SE  (.I(io_in[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[3]_SE  (.I(io_in[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[35]_SE  (.I(io_in[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[34]_SE  (.I(io_in[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[4]_SE  (.I(io_in[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[5]_SE  (.I(io_in[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[33]_SE  (.I(io_in[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[2]_SE  (.I(io_in[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[37]_SE  (.I(io_in[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[38]_SE  (.I(io_in[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[39]_SE  (.I(io_in[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[0]_SE  (.I(io_in[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[1]_SE  (.I(io_in[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[9]_SE  (.I(io_in[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[36]_SE  (.I(io_in[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[8]_SE  (.I(io_in[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[7]_SE  (.I(io_in[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[53]_SE  (.I(io_in[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[50]_SE  (.I(io_in[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[49]_SE  (.I(io_in[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[51]_SE  (.I(io_in[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[48]_SE  (.I(io_in[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[47]_SE  (.I(io_in[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[46]_SE  (.I(io_in[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[45]_SE  (.I(io_in[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[44]_SE  (.I(io_in[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[52]_SE  (.I(io_in[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[42]_SE  (.I(io_in[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[43]_SE  (.I(io_in[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[40]_SE  (.I(io_in[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[41]_SE  (.I(io_in[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[56]_SE  (.I(io_in[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[55]_SE  (.I(io_in[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[64]_SE  (.I(io_in[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[63]_SE  (.I(io_in[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[62]_SE  (.I(io_in[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[61]_SE  (.I(io_in[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[60]_SE  (.I(io_in[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[59]_SE  (.I(io_in[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[58]_SE  (.I(io_in[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[57]_SE  (.I(io_in[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[68]_SE  (.I(io_in[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[67]_SE  (.I(io_in[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[69]_SE  (.I(io_in[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[66]_SE  (.I(io_in[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[65]_SE  (.I(io_in[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[54]_SE  (.I(io_in[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[13]_SE  (.I(io_in[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[12]_SE  (.I(io_in[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[11]_SE  (.I(io_in[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[10]_SE  (.I(io_in[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[28]_SE  (.I(io_in[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[29]_SE  (.I(io_in[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[30]_SE  (.I(io_in[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[6]_SE  (.I(io_in[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09817__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09620__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09819__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09818__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09621__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09622__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09822__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09820__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09623__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09725__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09724__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09914__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09913__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09726__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09916__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09915__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09728__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09918__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09821__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09917__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09625__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09624__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09729__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09727__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09979__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09978__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09977__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10796__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10795__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10794__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10365__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10364__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10363__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10799__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09982__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10368__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10604__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10595__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10596__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10599__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10603__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10606__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10598__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10355__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10357__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10356__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10607__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10360__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10074__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09988__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09986__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10076__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10075__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10359__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09981__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09987__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10797__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10366__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10367__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10798__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10358__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09980__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09898__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09883__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09875__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09899__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09891__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09627__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09890__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09882__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09874__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09824__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09919__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09626__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09731__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09895__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09903__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09730__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09884__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09876__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09892__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09943__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09927__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09931__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09939__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09923__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09900__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10792__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09924__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09922__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09940__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09932__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09935__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10789__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10788__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10793__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10790__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10787__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09885__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09877__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09938__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09930__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09925__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09941__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09933__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09928__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09944__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09936__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09901__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09920__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09887__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09879__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09880__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09888__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09896__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09823__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09893__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09954__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09886__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10801__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10370__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09902__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09894__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09878__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09984__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10369__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09983__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10800__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09904__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10610__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10602__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10609__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10601__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09967__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09962__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09951__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09959__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09946__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09966__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09950__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09958__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10362__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10361__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10786__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10791__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09865__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09921__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09871__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09937__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09929__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09942__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09889__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09897__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09873__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09881__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09934__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09926__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09964__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09949__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09948__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09957__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09956__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09867__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09870__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09965__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09869__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09868__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09866__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09872__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10170__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10078__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10077__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10171__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10172__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10028__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10026__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10027__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10174__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10422__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10421__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10423__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10030__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10173__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10029__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09989__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10892__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10896__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10895__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10893__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09615__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09612__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09616__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09613__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10894__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10597__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09614__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10169__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09617__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10897__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10025__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10605__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10949__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10950__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10936__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10667__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10938__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10939__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10952__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10951__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10937__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10940__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10953__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10948__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10935__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10474__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10491__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10490__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10428__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10666__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10427__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10426__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10425__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10668__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10429__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10669__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10424__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10674__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10680__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10681__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10678__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10420__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10419__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09985__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10073__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10608__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10600__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09990__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10489__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10488__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09975__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09974__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09970__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10898__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10079__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09960__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10899__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09619__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09947__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09955__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09618__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10176__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09971__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09952__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09991__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09968__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09973__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09972__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09602__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09603__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09911__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09953__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09912__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09600__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09909__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09961__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09969__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09601__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09598__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09906__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09751__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09752__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09963__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10031__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09992__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10032__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09976__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10175__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10080__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09945__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09905__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09749__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09741__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09744__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09743__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09995__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10000__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10943__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10942__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10230__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09999__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10945__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10245__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10243__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10244__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10229__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10228__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09996__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09997__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10934__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10947__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10015__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10473__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10242__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10241__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10227__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10226__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10225__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10071__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10007__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10240__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09993__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09994__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10016__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10008__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10072__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10954__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09747__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09738__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09739__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09750__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09742__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09908__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09740__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09748__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09998__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09910__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09907__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09775__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09776__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10924__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10159__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10168__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10013__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10021__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10167__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10005__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10160__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10069__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10867__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10875__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10883__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10891__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10890__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10882__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10874__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10866__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10878__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10886__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10881__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10889__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10870__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10865__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10873__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10862__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10871__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10884__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10860__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10876__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10872__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10868__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10864__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10887__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10879__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10880__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10877__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10885__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10869__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10861__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10863__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10821__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10808__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10824__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10840__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10805__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10837__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10781__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10825__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10841__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10809__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10785__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10784__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10820__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10804__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10836__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10780__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10782__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10822__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10819__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10779__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10778__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10818__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10803__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10802__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10835__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10834__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10658__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10665__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10549__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10545__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10544__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10503__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10550__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10508__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10509__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10551__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10502__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10664__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10888__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10547__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10546__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10505__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10659__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10660__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10548__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10506__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10504__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10663__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10662__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10661__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10507__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10693__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10911__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10685__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10701__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10683__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10699__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10691__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10909__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10696__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10914__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10913__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10695__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10688__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10704__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10687__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10703__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10915__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10698__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10689__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10700__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10694__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10705__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10697__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10702__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10692__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10686__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10690__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10807__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10783__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10839__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10823__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10768__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10833__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10767__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10832__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10769__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10593__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10592__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10591__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10806__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10838__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10831__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10816__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10817__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10815__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10810__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10765__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10589__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10829__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10813__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10736__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10735__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10733__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10752__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10751__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10749__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10744__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10743__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10741__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10742__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10750__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10734__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10828__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10812__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10588__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10738__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10753__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10745__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10710__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10739__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10711__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10654__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10906__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10709__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10712__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10740__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10737__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10827__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10826__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10830__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10814__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10590__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10586__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10763__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10587__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10762__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10766__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10811__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10651__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10904__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10903__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10905__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10719__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10627__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10628__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10629__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10630__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10717__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10720__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10718__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10764__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10929__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10926__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10932__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10931__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10930__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09609__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09586__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09585__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09611__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10184__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10925__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10927__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10183__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10182__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09597__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09596__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10912__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10760__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09578__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09608__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09584__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10910__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10761__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10759__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09579__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09577__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10682__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10908__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10684__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09575__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10757__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09588__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09594__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09581__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10754__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09574__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10756__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09605__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10181__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09572__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09634__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09593__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09633__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09595__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09580__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10178__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09582__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09606__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09604__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09607__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09745__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09737__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10179__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10177__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09583__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09599__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09746__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09826__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10774__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10050__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09591__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10638__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10635__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10634__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10632__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09590__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09628__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09630__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09631__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10301__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10305__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10614__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10299__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10646__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10642__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10617__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10061__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10058__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10054__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10062__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10775__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10771__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10053__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10643__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10640__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10611__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10055__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10063__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10613__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10928__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10180__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09587__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09610__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10716__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10902__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10748__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10731__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10713__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10708__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10732__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10746__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10730__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10747__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10923__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09632__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10284__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10292__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10758__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10755__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09592__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09573__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10706__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10293__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10285__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09576__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10707__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09635__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10655__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10652__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10631__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10625__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10901__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10900__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10715__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10714__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10907__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10721__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10653__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10920__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10919__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10921__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10649__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10291__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10290__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10289__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10283__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10282__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10281__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10650__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10648__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10626__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10624__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10633__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10641__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10639__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10844__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09589__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09629__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10922__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10849__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10848__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10618__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10647__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10644__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10616__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10615__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10612__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10637__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10843__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10286__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10918__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10280__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10847__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10846__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10287__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10279__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10845__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10278__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10916__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10917__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10288__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10372__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10376__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10377__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10842__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10467__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10468__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10444__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10393__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10449__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10448__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10463__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10388__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10392__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10387__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10462__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10443__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10636__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10645__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10676__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10679__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10434__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10433__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10432__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10431__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10430__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10670__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10675__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10672__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10671__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10673__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10480__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10479__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10619__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10452__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10858__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10453__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10487__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10454__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10476__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10620__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10475__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10471__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10492__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10295__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10418__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10677__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10478__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10477__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10411__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10436__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10437__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10438__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10440__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10439__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10417__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10416__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10415__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10435__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10594__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10482__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10456__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10656__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10458__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10457__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10451__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10486__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10483__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10455__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10485__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10484__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10481__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10623__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10014__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10022__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10941__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10239__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10023__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10024__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10472__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10068__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10070__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10006__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10621__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10622__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10010__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10019__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10011__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10157__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09773__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10020__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10012__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10004__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10165__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10164__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10156__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09772__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09769__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10001__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10166__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10153__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10158__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10161__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09774__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10956__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10066__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10067__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10002__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10955__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10003__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10009__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10017__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10065__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10853__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10127__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10851__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09735__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09734__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09733__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09736__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10470__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10460__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10459__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10018__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10461__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10148__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10855__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10850__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10946__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09723__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09683__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09718__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10143__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10154__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10155__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10162__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10163__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09770__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09771__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10135__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09717__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09677__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09701__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10106__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10128__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10124__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10132__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10140__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10852__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10151__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10854__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10136__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10112__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10107__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09678__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09707__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09702__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10144__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10541__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10298__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10296__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10294__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10510__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10270__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10552__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10540__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10585__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10276__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10272__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10271__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10273__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10553__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10933__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10511__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10554__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10558__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10513__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10514__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10557__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10556__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10555__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10657__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10442__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10441__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10412__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10413__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10414__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10542__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10543__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10583__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10575__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10573__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10574__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10525__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10524__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10576__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10569__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10568__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10572__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10571__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10570__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10584__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10539__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10538__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10529__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10520__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10564__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10519__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10518__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10521__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10516__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10561__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10560__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10559__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10515__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10565__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10566__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10567__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10563__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10517__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10562__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10512__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10528__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10527__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10526__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10523__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10522__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10859__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10493__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10149__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10142__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10141__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10150__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10856__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09732__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10857__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10126__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10125__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10133__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10134__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10944__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10275__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10138__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10139__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10537__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10582__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10581__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10274__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10297__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10122__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10130__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10131__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10123__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10277__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10087__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09704__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09722__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09721__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09682__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09681__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09706__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09705__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10110__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10111__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09720__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09680__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10109__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10152__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10137__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10116__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10100__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09780__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10119__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10088__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10120__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10104__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09784__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09783__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10103__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10129__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10121__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10084__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09849__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10085__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09778__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09779__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10115__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10086__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10098__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10083__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10145__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10081__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09777__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10082__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10113__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10097__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09843__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09851__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09859__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09782__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09781__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10118__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10114__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10102__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10101__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10117__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09835__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10531__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10579__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10578__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10577__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10532__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10534__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10533__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10580__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10099__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10535__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10146__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10147__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10536__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10530__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10059__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10770__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10049__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09827__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10772__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10051__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10060__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10052__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10773__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10189__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10188__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10191__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10192__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09829__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09830__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10057__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10725__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09638__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10722__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10723__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10724__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10727__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09641__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09639__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09637__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09636__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09825__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09828__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10185__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10190__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10339__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10777__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10056__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10064__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10302__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09761__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09766__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09767__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10323__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10776__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09831__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10399__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09763__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09642__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09643__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10726__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10729__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10728__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09764__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09765__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09640__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09762__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10395__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10343__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10327__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09832__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09786__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09785__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09804__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09788__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09790__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09787__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10187__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10186__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10267__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10094__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09703__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10108__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09719__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09679__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10246__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10091__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10397__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09805__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09808__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09807__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09791__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10253__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10095__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10252__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10325__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09792__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09789__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09768__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10093__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10268__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10269__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10247__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09806__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09801__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09802__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09803__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10259__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10089__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10090__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10248__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10251__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10096__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10261__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10092__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10249__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10250__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10389__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10306__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10304__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10303__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10300__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10344__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10328__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10345__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10329__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10371__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10342__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10401__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10400__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10341__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10237__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10238__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10347__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10232__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10386__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10379__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10231__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10381__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10233__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10380__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10236__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10235__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10350__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10348__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10383__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10352__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10384__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10382__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10447__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10373__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10375__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10374__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10450__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10378__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10391__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10466__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10465__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10446__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10390__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10394__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10469__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10464__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10445__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10385__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10346__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10340__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10398__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10326__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10353__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10234__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10315__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10322__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10354__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10338__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10396__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10402__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10330__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10324__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10313__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10321__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10337__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10494__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10403__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10500__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10409__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10410__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10336__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10349__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10351__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10331__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10333__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10332__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10311__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10319__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10312__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10335__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10334__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10309__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10317__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10408__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10320__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10496__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10310__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10497__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10495__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10406__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10404__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10499__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10407__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10498__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10318__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10405__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10308__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10316__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10307__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10501__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10314__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10260__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09815__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10262__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09834__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09700__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09676__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09716__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10105__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09799__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09847__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09839__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09863__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09855__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09842__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10254__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10036__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09793__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09809__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10035__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09811__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09795__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09796__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09812__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10043__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10039__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09850__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09858__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10044__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09844__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09852__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09836__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10047__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10256__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10265__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10264__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10266__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10263__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10255__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09693__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09645__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09650__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09698__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10258__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10257__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09675__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10048__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09647__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09754__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09685__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09759__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09651__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09699__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09800__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09816__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09760__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09691__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09644__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09690__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10041__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10033__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09857__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09833__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09841__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09860__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09810__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09794__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09814__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09798__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10046__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10042__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10034__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09837__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09845__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09861__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09853__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09848__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10038__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09840__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09856__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09864__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09862__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09846__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09854__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09838__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09696__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09649__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09648__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10040__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09646__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09694__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10045__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09695__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09756__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09813__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09753__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09797__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09687__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09692__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09684__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09697__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09686__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09755__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09688__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09689__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09757__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09758__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10037__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09661__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09659__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10200__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09709__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10208__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09674__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09666__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09714__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09658__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09653__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10207__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10199__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10215__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10223__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09652__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09711__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09708__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09663__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09660__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10201__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10193__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10209__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09671__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10216__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09669__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09667__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09715__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09655__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10224__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10202__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10210__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10222__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10194__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10204__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10196__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10206__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10198__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10212__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10220__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10214__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10221__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10213__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10219__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10211__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10197__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10195__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10203__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10218__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10205__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09673__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09656__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09657__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09712__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09665__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09664__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09672__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09713__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09668__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09662__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09670__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09654__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09710__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10217__CLK (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[2]_D  (.I(\u_arbiter.i_wb_cpu_ack ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08921__A1 (.I(\u_arbiter.i_wb_cpu_ack ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08197__A1 (.I(\u_arbiter.i_wb_cpu_ack ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08012__A1 (.I(\u_arbiter.i_wb_cpu_ack ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06485__A1 (.I(\u_arbiter.i_wb_cpu_ack ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06469__A1 (.I(\u_arbiter.i_wb_cpu_ack ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08607__I1 (.I(\u_arbiter.i_wb_cpu_dbus_adr[23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08605__I0 (.I(\u_arbiter.i_wb_cpu_dbus_adr[23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05013__A1 (.I(\u_arbiter.i_wb_cpu_dbus_adr[23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08611__I1 (.I(\u_arbiter.i_wb_cpu_dbus_adr[25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08609__I0 (.I(\u_arbiter.i_wb_cpu_dbus_adr[25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05020__A1 (.I(\u_arbiter.i_wb_cpu_dbus_adr[25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08619__I1 (.I(\u_arbiter.i_wb_cpu_dbus_adr[29] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08617__I0 (.I(\u_arbiter.i_wb_cpu_dbus_adr[29] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05036__A1 (.I(\u_arbiter.i_wb_cpu_dbus_adr[29] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08568__I1 (.I(\u_arbiter.i_wb_cpu_dbus_adr[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08566__I0 (.I(\u_arbiter.i_wb_cpu_dbus_adr[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04930__A1 (.I(\u_arbiter.i_wb_cpu_dbus_adr[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[6]_SI  (.I(\u_arbiter.i_wb_cpu_dbus_dat[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08025__A1 (.I(\u_arbiter.i_wb_cpu_dbus_dat[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08018__A1 (.I(\u_arbiter.i_wb_cpu_dbus_dat[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08015__B2 (.I(\u_arbiter.i_wb_cpu_dbus_dat[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08009__A1 (.I(\u_arbiter.i_wb_cpu_dbus_dat[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06479__A1 (.I(\u_arbiter.i_wb_cpu_dbus_dat[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05904__I0 (.I(\u_arbiter.i_wb_cpu_dbus_dat[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[20]_SI  (.I(\u_arbiter.i_wb_cpu_dbus_dat[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08072__B2 (.I(\u_arbiter.i_wb_cpu_dbus_dat[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08069__A1 (.I(\u_arbiter.i_wb_cpu_dbus_dat[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[22]_SI  (.I(\u_arbiter.i_wb_cpu_dbus_dat[16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08078__B2 (.I(\u_arbiter.i_wb_cpu_dbus_dat[16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08074__A1 (.I(\u_arbiter.i_wb_cpu_dbus_dat[16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05904__I2 (.I(\u_arbiter.i_wb_cpu_dbus_dat[16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[7]_SI  (.I(\u_arbiter.i_wb_cpu_dbus_dat[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08025__A2 (.I(\u_arbiter.i_wb_cpu_dbus_dat[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08020__A1 (.I(\u_arbiter.i_wb_cpu_dbus_dat[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08018__A2 (.I(\u_arbiter.i_wb_cpu_dbus_dat[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08011__A1 (.I(\u_arbiter.i_wb_cpu_dbus_dat[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06479__A2 (.I(\u_arbiter.i_wb_cpu_dbus_dat[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[30]_SI  (.I(\u_arbiter.i_wb_cpu_dbus_dat[24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08100__A1 (.I(\u_arbiter.i_wb_cpu_dbus_dat[24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08096__A1 (.I(\u_arbiter.i_wb_cpu_dbus_dat[24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05904__I3 (.I(\u_arbiter.i_wb_cpu_dbus_dat[24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[8]_SI  (.I(\u_arbiter.i_wb_cpu_dbus_dat[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08027__A1 (.I(\u_arbiter.i_wb_cpu_dbus_dat[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08025__A3 (.I(\u_arbiter.i_wb_cpu_dbus_dat[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08017__A1 (.I(\u_arbiter.i_wb_cpu_dbus_dat[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06479__A3 (.I(\u_arbiter.i_wb_cpu_dbus_dat[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[11]_SI  (.I(\u_arbiter.i_wb_cpu_dbus_dat[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08046__A1 (.I(\u_arbiter.i_wb_cpu_dbus_dat[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08041__A1 (.I(\u_arbiter.i_wb_cpu_dbus_dat[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06481__A1 (.I(\u_arbiter.i_wb_cpu_dbus_dat[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05886__A1 (.I(\u_arbiter.i_wb_cpu_dbus_dat[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[12]_SI  (.I(\u_arbiter.i_wb_cpu_dbus_dat[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08048__B2 (.I(\u_arbiter.i_wb_cpu_dbus_dat[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06475__A1 (.I(\u_arbiter.i_wb_cpu_dbus_dat[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[14]_SI  (.I(\u_arbiter.i_wb_cpu_dbus_dat[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08055__B2 (.I(\u_arbiter.i_wb_cpu_dbus_dat[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08051__A1 (.I(\u_arbiter.i_wb_cpu_dbus_dat[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05904__I1 (.I(\u_arbiter.i_wb_cpu_dbus_dat[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08658__A1 (.I(\u_arbiter.i_wb_cpu_ibus_adr[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05987__A1 (.I(\u_arbiter.i_wb_cpu_ibus_adr[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05982__A1 (.I(\u_arbiter.i_wb_cpu_ibus_adr[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05921__A1 (.I(\u_arbiter.i_wb_cpu_ibus_adr[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05898__A1 (.I(\u_arbiter.i_wb_cpu_ibus_adr[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05867__A1 (.I(\u_arbiter.i_wb_cpu_ibus_adr[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04908__A1 (.I(\u_arbiter.i_wb_cpu_ibus_adr[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08660__A1 (.I(\u_arbiter.i_wb_cpu_ibus_adr[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08658__B2 (.I(\u_arbiter.i_wb_cpu_ibus_adr[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08196__A2 (.I(\u_arbiter.i_wb_cpu_ibus_adr[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06470__A2 (.I(\u_arbiter.i_wb_cpu_ibus_adr[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04910__A1 (.I(\u_arbiter.i_wb_cpu_ibus_adr[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[3]_D  (.I(\u_arbiter.i_wb_cpu_rdt[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08474__I1 (.I(\u_arbiter.i_wb_cpu_rdt[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08172__I0 (.I(\u_arbiter.i_wb_cpu_rdt[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08154__A2 (.I(\u_arbiter.i_wb_cpu_rdt[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08015__A1 (.I(\u_arbiter.i_wb_cpu_rdt[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[13]_D  (.I(\u_arbiter.i_wb_cpu_rdt[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08307__I1 (.I(\u_arbiter.i_wb_cpu_rdt[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08142__I0 (.I(\u_arbiter.i_wb_cpu_rdt[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08061__A1 (.I(\u_arbiter.i_wb_cpu_rdt[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[14]_D  (.I(\u_arbiter.i_wb_cpu_rdt[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08390__I1 (.I(\u_arbiter.i_wb_cpu_rdt[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08141__I0 (.I(\u_arbiter.i_wb_cpu_rdt[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08064__A1 (.I(\u_arbiter.i_wb_cpu_rdt[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[15]_D  (.I(\u_arbiter.i_wb_cpu_rdt[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08395__A2 (.I(\u_arbiter.i_wb_cpu_rdt[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08235__I0 (.I(\u_arbiter.i_wb_cpu_rdt[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08151__A2 (.I(\u_arbiter.i_wb_cpu_rdt[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08067__A1 (.I(\u_arbiter.i_wb_cpu_rdt[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[16]_D  (.I(\u_arbiter.i_wb_cpu_rdt[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08407__A2 (.I(\u_arbiter.i_wb_cpu_rdt[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08203__I0 (.I(\u_arbiter.i_wb_cpu_rdt[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08185__A2 (.I(\u_arbiter.i_wb_cpu_rdt[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08070__A1 (.I(\u_arbiter.i_wb_cpu_rdt[13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[17]_D  (.I(\u_arbiter.i_wb_cpu_rdt[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08415__I1 (.I(\u_arbiter.i_wb_cpu_rdt[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08175__I0 (.I(\u_arbiter.i_wb_cpu_rdt[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08167__A2 (.I(\u_arbiter.i_wb_cpu_rdt[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08072__A1 (.I(\u_arbiter.i_wb_cpu_rdt[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[18]_D  (.I(\u_arbiter.i_wb_cpu_rdt[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08519__I1 (.I(\u_arbiter.i_wb_cpu_rdt[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08178__A2 (.I(\u_arbiter.i_wb_cpu_rdt[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08168__I0 (.I(\u_arbiter.i_wb_cpu_rdt[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08075__A1 (.I(\u_arbiter.i_wb_cpu_rdt[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[19]_D  (.I(\u_arbiter.i_wb_cpu_rdt[16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08943__I0 (.I(\u_arbiter.i_wb_cpu_rdt[16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08474__I0 (.I(\u_arbiter.i_wb_cpu_rdt[16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08078__A1 (.I(\u_arbiter.i_wb_cpu_rdt[16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[20]_D  (.I(\u_arbiter.i_wb_cpu_rdt[17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08945__I0 (.I(\u_arbiter.i_wb_cpu_rdt[17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08488__I0 (.I(\u_arbiter.i_wb_cpu_rdt[17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08080__A1 (.I(\u_arbiter.i_wb_cpu_rdt[17] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[21]_D  (.I(\u_arbiter.i_wb_cpu_rdt[18] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08947__I0 (.I(\u_arbiter.i_wb_cpu_rdt[18] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08498__I0 (.I(\u_arbiter.i_wb_cpu_rdt[18] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08083__A1 (.I(\u_arbiter.i_wb_cpu_rdt[18] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[4]_D  (.I(\u_arbiter.i_wb_cpu_rdt[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08488__I1 (.I(\u_arbiter.i_wb_cpu_rdt[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08201__A2 (.I(\u_arbiter.i_wb_cpu_rdt[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08155__I0 (.I(\u_arbiter.i_wb_cpu_rdt[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08022__A1 (.I(\u_arbiter.i_wb_cpu_rdt[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[23]_D  (.I(\u_arbiter.i_wb_cpu_rdt[20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08951__I0 (.I(\u_arbiter.i_wb_cpu_rdt[20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08254__I0 (.I(\u_arbiter.i_wb_cpu_rdt[20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08089__A1 (.I(\u_arbiter.i_wb_cpu_rdt[20] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[24]_D  (.I(\u_arbiter.i_wb_cpu_rdt[21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08953__I0 (.I(\u_arbiter.i_wb_cpu_rdt[21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08265__I0 (.I(\u_arbiter.i_wb_cpu_rdt[21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08091__A1 (.I(\u_arbiter.i_wb_cpu_rdt[21] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[25]_D  (.I(\u_arbiter.i_wb_cpu_rdt[22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08955__I0 (.I(\u_arbiter.i_wb_cpu_rdt[22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08277__I0 (.I(\u_arbiter.i_wb_cpu_rdt[22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08094__A1 (.I(\u_arbiter.i_wb_cpu_rdt[22] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[26]_D  (.I(\u_arbiter.i_wb_cpu_rdt[23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08957__I0 (.I(\u_arbiter.i_wb_cpu_rdt[23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08346__I0 (.I(\u_arbiter.i_wb_cpu_rdt[23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08097__A1 (.I(\u_arbiter.i_wb_cpu_rdt[23] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[27]_D  (.I(\u_arbiter.i_wb_cpu_rdt[24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08959__I0 (.I(\u_arbiter.i_wb_cpu_rdt[24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08359__I0 (.I(\u_arbiter.i_wb_cpu_rdt[24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08099__A1 (.I(\u_arbiter.i_wb_cpu_rdt[24] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[28]_D  (.I(\u_arbiter.i_wb_cpu_rdt[25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08961__I0 (.I(\u_arbiter.i_wb_cpu_rdt[25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08375__A2 (.I(\u_arbiter.i_wb_cpu_rdt[25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08104__A1 (.I(\u_arbiter.i_wb_cpu_rdt[25] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[29]_D  (.I(\u_arbiter.i_wb_cpu_rdt[26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08963__I0 (.I(\u_arbiter.i_wb_cpu_rdt[26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08307__I0 (.I(\u_arbiter.i_wb_cpu_rdt[26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08106__A1 (.I(\u_arbiter.i_wb_cpu_rdt[26] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[30]_D  (.I(\u_arbiter.i_wb_cpu_rdt[27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08965__I0 (.I(\u_arbiter.i_wb_cpu_rdt[27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08390__I0 (.I(\u_arbiter.i_wb_cpu_rdt[27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08109__A1 (.I(\u_arbiter.i_wb_cpu_rdt[27] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[31]_D  (.I(\u_arbiter.i_wb_cpu_rdt[28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08967__I0 (.I(\u_arbiter.i_wb_cpu_rdt[28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08396__A2 (.I(\u_arbiter.i_wb_cpu_rdt[28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08112__A1 (.I(\u_arbiter.i_wb_cpu_rdt[28] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[32]_D  (.I(\u_arbiter.i_wb_cpu_rdt[29] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08969__I0 (.I(\u_arbiter.i_wb_cpu_rdt[29] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08408__A2 (.I(\u_arbiter.i_wb_cpu_rdt[29] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08115__A1 (.I(\u_arbiter.i_wb_cpu_rdt[29] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[5]_D  (.I(\u_arbiter.i_wb_cpu_rdt[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08498__I1 (.I(\u_arbiter.i_wb_cpu_rdt[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08163__I0 (.I(\u_arbiter.i_wb_cpu_rdt[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08029__A1 (.I(\u_arbiter.i_wb_cpu_rdt[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[33]_D  (.I(\u_arbiter.i_wb_cpu_rdt[30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08971__I0 (.I(\u_arbiter.i_wb_cpu_rdt[30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08415__I0 (.I(\u_arbiter.i_wb_cpu_rdt[30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08118__A1 (.I(\u_arbiter.i_wb_cpu_rdt[30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[34]_D  (.I(\u_arbiter.i_wb_cpu_rdt[31] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08973__I0 (.I(\u_arbiter.i_wb_cpu_rdt[31] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08519__I0 (.I(\u_arbiter.i_wb_cpu_rdt[31] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08120__A1 (.I(\u_arbiter.i_wb_cpu_rdt[31] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[7]_D  (.I(\u_arbiter.i_wb_cpu_rdt[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08254__I1 (.I(\u_arbiter.i_wb_cpu_rdt[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08162__I0 (.I(\u_arbiter.i_wb_cpu_rdt[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08043__A1 (.I(\u_arbiter.i_wb_cpu_rdt[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[8]_D  (.I(\u_arbiter.i_wb_cpu_rdt[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08309__I0 (.I(\u_arbiter.i_wb_cpu_rdt[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08265__I1 (.I(\u_arbiter.i_wb_cpu_rdt[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08159__A2 (.I(\u_arbiter.i_wb_cpu_rdt[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08045__A1 (.I(\u_arbiter.i_wb_cpu_rdt[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[9]_D  (.I(\u_arbiter.i_wb_cpu_rdt[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08277__I1 (.I(\u_arbiter.i_wb_cpu_rdt[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08156__I0 (.I(\u_arbiter.i_wb_cpu_rdt[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08048__A1 (.I(\u_arbiter.i_wb_cpu_rdt[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[10]_D  (.I(\u_arbiter.i_wb_cpu_rdt[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08430__A2 (.I(\u_arbiter.i_wb_cpu_rdt[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08346__I1 (.I(\u_arbiter.i_wb_cpu_rdt[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08144__I0 (.I(\u_arbiter.i_wb_cpu_rdt[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08052__A1 (.I(\u_arbiter.i_wb_cpu_rdt[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[11]_D  (.I(\u_arbiter.i_wb_cpu_rdt[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08359__I1 (.I(\u_arbiter.i_wb_cpu_rdt[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08188__I0 (.I(\u_arbiter.i_wb_cpu_rdt[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08147__A2 (.I(\u_arbiter.i_wb_cpu_rdt[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08055__A1 (.I(\u_arbiter.i_wb_cpu_rdt[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[12]_D  (.I(\u_arbiter.i_wb_cpu_rdt[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08401__A2 (.I(\u_arbiter.i_wb_cpu_rdt[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08376__A2 (.I(\u_arbiter.i_wb_cpu_rdt[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08143__I0 (.I(\u_arbiter.i_wb_cpu_rdt[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08058__A1 (.I(\u_arbiter.i_wb_cpu_rdt[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[54]_SI  (.I(\u_arbiter.o_wb_cpu_adr[16] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[68]_SI  (.I(\u_arbiter.o_wb_cpu_adr[30] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[69]_SI  (.I(\u_arbiter.o_wb_cpu_adr[31] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05825__I (.I(\u_cpu.cpu.alu.i_rs1 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05995__A2 (.I(\u_cpu.cpu.bne_or_bge ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05871__A1 (.I(\u_cpu.cpu.bne_or_bge ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05850__I (.I(\u_cpu.cpu.bne_or_bge ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04883__A2 (.I(\u_cpu.cpu.bne_or_bge ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04857__A4 (.I(\u_cpu.cpu.bne_or_bge ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04845__A3 (.I(\u_cpu.cpu.bne_or_bge ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08919__A1 (.I(\u_cpu.cpu.bufreg.i_sh_signed ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08624__A1 (.I(\u_cpu.cpu.bufreg.i_sh_signed ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05824__A2 (.I(\u_cpu.cpu.bufreg.i_sh_signed ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08005__C (.I(\u_cpu.cpu.bufreg.lsb[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05997__A1 (.I(\u_cpu.cpu.bufreg.lsb[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05995__A1 (.I(\u_cpu.cpu.bufreg.lsb[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05904__S0 (.I(\u_cpu.cpu.bufreg.lsb[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05879__I (.I(\u_cpu.cpu.bufreg.lsb[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04842__A1 (.I(\u_cpu.cpu.bufreg.lsb[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08630__A1 (.I(\u_cpu.cpu.bufreg.lsb[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08006__A1 (.I(\u_cpu.cpu.bufreg.lsb[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08005__A1 (.I(\u_cpu.cpu.bufreg.lsb[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05996__A1 (.I(\u_cpu.cpu.bufreg.lsb[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05964__I (.I(\u_cpu.cpu.bufreg.lsb[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05904__S1 (.I(\u_cpu.cpu.bufreg.lsb[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04842__A2 (.I(\u_cpu.cpu.bufreg.lsb[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09395__A1 (.I(\u_cpu.cpu.ctrl.i_iscomp ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05896__A2 (.I(\u_cpu.cpu.ctrl.i_iscomp ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05895__A2 (.I(\u_cpu.cpu.ctrl.i_iscomp ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08686__A1 (.I(\u_cpu.cpu.ctrl.o_ibus_adr[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08684__B2 (.I(\u_cpu.cpu.ctrl.o_ibus_adr[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04978__A2 (.I(\u_cpu.cpu.ctrl.o_ibus_adr[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04977__A1 (.I(\u_cpu.cpu.ctrl.o_ibus_adr[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04975__A1 (.I(\u_cpu.cpu.ctrl.o_ibus_adr[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04974__A1 (.I(\u_cpu.cpu.ctrl.o_ibus_adr[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08689__A1 (.I(\u_cpu.cpu.ctrl.o_ibus_adr[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08686__B2 (.I(\u_cpu.cpu.ctrl.o_ibus_adr[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04978__A1 (.I(\u_cpu.cpu.ctrl.o_ibus_adr[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04977__B (.I(\u_cpu.cpu.ctrl.o_ibus_adr[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09386__A1 (.I(\u_cpu.cpu.decode.co_ebreak ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05861__A2 (.I(\u_cpu.cpu.decode.co_ebreak ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04886__A2 (.I(\u_cpu.cpu.decode.co_ebreak ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04855__I (.I(\u_cpu.cpu.decode.co_ebreak ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05860__I (.I(\u_cpu.cpu.decode.op21 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04868__A1 (.I(\u_cpu.cpu.decode.op21 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04857__A3 (.I(\u_cpu.cpu.decode.op21 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04856__A1 (.I(\u_cpu.cpu.decode.op21 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04851__A1 (.I(\u_cpu.cpu.decode.op21 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08445__A2 (.I(\u_cpu.cpu.decode.opcode[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08424__B (.I(\u_cpu.cpu.decode.opcode[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08207__A1 (.I(\u_cpu.cpu.decode.opcode[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05975__A1 (.I(\u_cpu.cpu.decode.opcode[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05972__A2 (.I(\u_cpu.cpu.decode.opcode[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05919__A1 (.I(\u_cpu.cpu.decode.opcode[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05830__A2 (.I(\u_cpu.cpu.decode.opcode[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08961__I1 (.I(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08400__A2 (.I(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08143__I1 (.I(\u_cpu.cpu.genblk1.align.ibus_rdt_concat[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[1]_D  (.I(\u_cpu.cpu.genblk3.csr.i_mtip ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08524__A3 (.I(\u_cpu.cpu.genblk3.csr.i_mtip ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09397__A1 (.I(\u_cpu.cpu.genblk3.csr.o_new_irq ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09381__A1 (.I(\u_cpu.cpu.genblk3.csr.o_new_irq ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09373__B (.I(\u_cpu.cpu.genblk3.csr.o_new_irq ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09364__A1 (.I(\u_cpu.cpu.genblk3.csr.o_new_irq ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05983__A1 (.I(\u_cpu.cpu.genblk3.csr.o_new_irq ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04867__A1 (.I(\u_cpu.cpu.genblk3.csr.o_new_irq ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04858__I (.I(\u_cpu.cpu.genblk3.csr.o_new_irq ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08824__A1 (.I(\u_cpu.cpu.immdec.imm11_7[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08811__I1 (.I(\u_cpu.cpu.immdec.imm11_7[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08729__A1 (.I(\u_cpu.cpu.immdec.imm11_7[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06330__A1 (.I(\u_cpu.cpu.immdec.imm11_7[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06254__A1 (.I(\u_cpu.cpu.immdec.imm11_7[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06013__A1 (.I(\u_cpu.cpu.immdec.imm11_7[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05991__A2 (.I(\u_cpu.cpu.immdec.imm11_7[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08829__A1 (.I(\u_cpu.cpu.immdec.imm11_7[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08820__A1 (.I(\u_cpu.cpu.immdec.imm11_7[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06330__A2 (.I(\u_cpu.cpu.immdec.imm11_7[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06157__A1 (.I(\u_cpu.cpu.immdec.imm11_7[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06078__A1 (.I(\u_cpu.cpu.immdec.imm11_7[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06017__A1 (.I(\u_cpu.cpu.immdec.imm11_7[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05991__A3 (.I(\u_cpu.cpu.immdec.imm11_7[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08486__A1 (.I(\u_cpu.cpu.immdec.imm19_12_20[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08472__A1 (.I(\u_cpu.cpu.immdec.imm19_12_20[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04881__A1 (.I(\u_cpu.cpu.immdec.imm19_12_20[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08513__A2 (.I(\u_cpu.cpu.immdec.imm24_20[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08338__A1 (.I(\u_cpu.cpu.immdec.imm24_20[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05832__B (.I(\u_cpu.cpu.immdec.imm24_20[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04863__A1 (.I(\u_cpu.cpu.immdec.imm24_20[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08341__A1 (.I(\u_cpu.cpu.immdec.imm24_20[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08337__A1 (.I(\u_cpu.cpu.immdec.imm24_20[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04888__A1 (.I(\u_cpu.cpu.immdec.imm24_20[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08363__A1 (.I(\u_cpu.cpu.immdec.imm24_20[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08355__A1 (.I(\u_cpu.cpu.immdec.imm24_20[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04875__A1 (.I(\u_cpu.cpu.immdec.imm24_20[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08837__A1 (.I(\u_cpu.cpu.immdec.imm30_25[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08380__A1 (.I(\u_cpu.cpu.immdec.imm30_25[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08363__B2 (.I(\u_cpu.cpu.immdec.imm30_25[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08520__A1 (.I(\u_cpu.cpu.immdec.imm31 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05911__A1 (.I(\u_cpu.cpu.immdec.imm31 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05834__A2 (.I(\u_cpu.cpu.immdec.imm31 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09386__A3 (.I(\u_cpu.cpu.mem_bytecnt[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08005__B (.I(\u_cpu.cpu.mem_bytecnt[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07679__A1 (.I(\u_cpu.cpu.mem_bytecnt[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07678__A1 (.I(\u_cpu.cpu.mem_bytecnt[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07677__A1 (.I(\u_cpu.cpu.mem_bytecnt[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05914__A2 (.I(\u_cpu.cpu.mem_bytecnt[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05903__B1 (.I(\u_cpu.cpu.mem_bytecnt[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05855__A3 (.I(\u_cpu.cpu.mem_bytecnt[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09386__A2 (.I(\u_cpu.cpu.mem_bytecnt[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08006__A2 (.I(\u_cpu.cpu.mem_bytecnt[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08005__A2 (.I(\u_cpu.cpu.mem_bytecnt[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07743__A1 (.I(\u_cpu.cpu.mem_bytecnt[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07680__A1 (.I(\u_cpu.cpu.mem_bytecnt[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05916__A1 (.I(\u_cpu.cpu.mem_bytecnt[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05903__A2 (.I(\u_cpu.cpu.mem_bytecnt[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05855__A1 (.I(\u_cpu.cpu.mem_bytecnt[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10940__D (.I(\u_cpu.cpu.o_wdata0 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06188__I1 (.I(\u_cpu.cpu.o_wdata0 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06065__A2 (.I(\u_cpu.cpu.o_wdata0 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10954__D (.I(\u_cpu.cpu.o_wdata1 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07729__A1 (.I(\u_cpu.cpu.state.genblk1.misalign_trap_sync_r ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06472__A1 (.I(\u_cpu.cpu.state.genblk1.misalign_trap_sync_r ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04867__A2 (.I(\u_cpu.cpu.state.genblk1.misalign_trap_sync_r ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04859__I (.I(\u_cpu.cpu.state.genblk1.misalign_trap_sync_r ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07745__A1 (.I(\u_cpu.cpu.state.init_done ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06487__A1 (.I(\u_cpu.cpu.state.init_done ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05983__A2 (.I(\u_cpu.cpu.state.init_done ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05968__A1 (.I(\u_cpu.cpu.state.init_done ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05888__A1 (.I(\u_cpu.cpu.state.init_done ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05880__A2 (.I(\u_cpu.cpu.state.init_done ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07683__A1 (.I(\u_cpu.cpu.state.o_cnt_r[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07675__A2 (.I(\u_cpu.cpu.state.o_cnt_r[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07674__A2 (.I(\u_cpu.cpu.state.o_cnt_r[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05966__A4 (.I(\u_cpu.cpu.state.o_cnt_r[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05857__A2 (.I(\u_cpu.cpu.state.o_cnt_r[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05820__A4 (.I(\u_cpu.cpu.state.o_cnt_r[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06558__A1 (.I(\u_cpu.rf_ram.memory[119][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05257__I3 (.I(\u_cpu.rf_ram.memory[119][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06562__A1 (.I(\u_cpu.rf_ram.memory[119][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05433__I3 (.I(\u_cpu.rf_ram.memory[119][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06566__A1 (.I(\u_cpu.rf_ram.memory[119][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05609__I3 (.I(\u_cpu.rf_ram.memory[119][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07837__A1 (.I(\u_cpu.rf_ram.memory[120][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05605__I0 (.I(\u_cpu.rf_ram.memory[120][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07515__A1 (.I(\u_cpu.rf_ram.memory[128][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05373__I0 (.I(\u_cpu.rf_ram.memory[128][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07521__A1 (.I(\u_cpu.rf_ram.memory[128][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05637__I0 (.I(\u_cpu.rf_ram.memory[128][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07486__A1 (.I(\u_cpu.rf_ram.memory[22][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05083__I2 (.I(\u_cpu.rf_ram.memory[22][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07489__A1 (.I(\u_cpu.rf_ram.memory[22][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05213__I2 (.I(\u_cpu.rf_ram.memory[22][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07498__A1 (.I(\u_cpu.rf_ram.memory[22][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05477__I2 (.I(\u_cpu.rf_ram.memory[22][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07501__A1 (.I(\u_cpu.rf_ram.memory[22][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05565__I2 (.I(\u_cpu.rf_ram.memory[22][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07504__A1 (.I(\u_cpu.rf_ram.memory[22][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05653__I2 (.I(\u_cpu.rf_ram.memory[22][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06792__A1 (.I(\u_cpu.rf_ram.memory[29][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05092__I1 (.I(\u_cpu.rf_ram.memory[29][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06798__A1 (.I(\u_cpu.rf_ram.memory[29][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05305__I1 (.I(\u_cpu.rf_ram.memory[29][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06801__A1 (.I(\u_cpu.rf_ram.memory[29][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05393__I1 (.I(\u_cpu.rf_ram.memory[29][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06804__A1 (.I(\u_cpu.rf_ram.memory[29][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05481__I1 (.I(\u_cpu.rf_ram.memory[29][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06807__A1 (.I(\u_cpu.rf_ram.memory[29][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05569__I1 (.I(\u_cpu.rf_ram.memory[29][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06810__A1 (.I(\u_cpu.rf_ram.memory[29][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05657__I1 (.I(\u_cpu.rf_ram.memory[29][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08648__A1 (.I(\u_cpu.rf_ram.memory[30][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05569__I2 (.I(\u_cpu.rf_ram.memory[30][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07290__A1 (.I(\u_cpu.rf_ram.memory[39][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05235__I3 (.I(\u_cpu.rf_ram.memory[39][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07292__A1 (.I(\u_cpu.rf_ram.memory[39][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05323__I3 (.I(\u_cpu.rf_ram.memory[39][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07294__A1 (.I(\u_cpu.rf_ram.memory[39][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05411__I3 (.I(\u_cpu.rf_ram.memory[39][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07300__A1 (.I(\u_cpu.rf_ram.memory[39][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05675__I3 (.I(\u_cpu.rf_ram.memory[39][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09223__A1 (.I(\u_cpu.rf_ram.memory[59][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05316__I3 (.I(\u_cpu.rf_ram.memory[59][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09229__A1 (.I(\u_cpu.rf_ram.memory[59][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05580__I3 (.I(\u_cpu.rf_ram.memory[59][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07751__A1 (.I(\u_cpu.rf_ram.memory[92][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05261__I0 (.I(\u_cpu.rf_ram.memory[92][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07753__A1 (.I(\u_cpu.rf_ram.memory[92][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05349__I0 (.I(\u_cpu.rf_ram.memory[92][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06021__I (.I(\u_cpu.rf_ram_if.genblk1.wtrig0_r ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06014__A1 (.I(\u_cpu.rf_ram_if.genblk1.wtrig0_r ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06003__I (.I(\u_cpu.rf_ram_if.genblk1.wtrig0_r ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06000__A1 (.I(\u_cpu.rf_ram_if.genblk1.wtrig0_r ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05999__B (.I(\u_cpu.rf_ram_if.genblk1.wtrig0_r ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10945__D (.I(\u_cpu.rf_ram_if.rtrig0 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09565__A3 (.I(\u_cpu.rf_ram_if.rtrig0 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06014__B1 (.I(\u_cpu.rf_ram_if.rtrig0 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04887__B (.I(\u_cpu.rf_ram_if.rtrig0 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04881__A2 (.I(\u_cpu.rf_ram_if.rtrig0 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04865__A2 (.I(\u_cpu.rf_ram_if.rtrig0 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__04862__A1 (.I(\u_cpu.rf_ram_if.rtrig0 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10952__D (.I(\u_cpu.rf_ram_if.wdata1_r[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06184__I1 (.I(\u_cpu.rf_ram_if.wdata1_r[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06058__A2 (.I(\u_cpu.rf_ram_if.wdata1_r[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[25]_CLK  (.I(\u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[24]_CLK  (.I(\u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[23]_CLK  (.I(\u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[22]_CLK  (.I(\u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[21]_CLK  (.I(\u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[20]_CLK  (.I(\u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[19]_CLK  (.I(\u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[18]_CLK  (.I(\u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[17]_CLK  (.I(\u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[16]_CLK  (.I(\u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[15]_CLK  (.I(\u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[14]_CLK  (.I(\u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[26]_CLK  (.I(\u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[32]_CLK  (.I(\u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[33]_CLK  (.I(\u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[28]_CLK  (.I(\u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[27]_CLK  (.I(\u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[29]_CLK  (.I(\u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[30]_CLK  (.I(\u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[31]_CLK  (.I(\u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[11]_CLK  (.I(\u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[12]_CLK  (.I(\u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[13]_CLK  (.I(\u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[10]_CLK  (.I(\u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[68]_CLK  (.I(\u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[67]_CLK  (.I(\u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[65]_CLK  (.I(\u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[66]_CLK  (.I(\u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[57]_CLK  (.I(\u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[56]_CLK  (.I(\u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[69]_CLK  (.I(\u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[64]_CLK  (.I(\u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.output_buffers[3]_I  (.I(\u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.out_flop_CLKN  (.I(\u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[61]_CLK  (.I(\u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[62]_CLK  (.I(\u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[63]_CLK  (.I(\u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[60]_CLK  (.I(\u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[59]_CLK  (.I(\u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[58]_CLK  (.I(\u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[40]_CLK  (.I(\u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[54]_CLK  (.I(\u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[45]_CLK  (.I(\u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[50]_CLK  (.I(\u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[49]_CLK  (.I(\u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[48]_CLK  (.I(\u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[47]_CLK  (.I(\u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[46]_CLK  (.I(\u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[51]_CLK  (.I(\u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[52]_CLK  (.I(\u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[53]_CLK  (.I(\u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[43]_CLK  (.I(\u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[44]_CLK  (.I(\u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[42]_CLK  (.I(\u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[41]_CLK  (.I(\u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[39]_CLK  (.I(\u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[38]_CLK  (.I(\u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[0]_CLK  (.I(\u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[1]_CLK  (.I(\u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[34]_CLK  (.I(\u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[35]_CLK  (.I(\u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[9]_CLK  (.I(\u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[37]_CLK  (.I(\u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[36]_CLK  (.I(\u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[6]_CLK  (.I(\u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[7]_CLK  (.I(\u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[8]_CLK  (.I(\u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[5]_CLK  (.I(\u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[4]_CLK  (.I(\u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[3]_CLK  (.I(\u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[2]_CLK  (.I(\u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[55]_CLK  (.I(\u_scanchain_local.clk ));
 gf180mcu_fd_sc_mcu7t5v0__antenna \ANTENNA_u_scanchain_local.scan_flop[42]_D  (.I(\u_scanchain_local.module_data_in[41] ));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_1_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_1_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_3_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_4_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_4_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_4_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_5_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_5_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_6_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_6_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_9_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_10_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_11_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_11_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_14_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_14_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_15_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_16_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_17_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_18_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_19_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_20_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_20_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_21_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_22_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_23_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_24_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_25_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_26_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_26_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_27_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_28_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_28_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_28_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_29_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_29_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_30_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_30_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_30_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_31_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_32_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_32_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_32_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_33_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_34_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_35_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_36_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_36_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_37_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_38_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_39_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_40_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_41_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_41_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_41_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_41_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_43_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_43_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_44_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_45_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_45_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_45_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_46_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_46_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_47_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_50_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_51_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_51_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_52_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_53_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_54_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_54_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_56_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_57_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_58_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_60_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_61_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_62_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_64_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_65_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_66_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_66_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_35 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_35 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_79_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_81_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_88_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_90_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_90_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_91_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_92_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_92_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_93_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_93_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_94_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_98_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_35 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_35 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_104_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_108_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_109_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_110_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_110_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_111_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_111_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_112_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_112_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_112_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_113_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_114_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_114_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_115_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_116_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_117_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_118_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_118_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_120_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_120_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_120_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_120_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_121_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_121_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_122_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_122_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_122_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_123_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_123_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_124_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_124_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_126_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_126_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_127_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_127_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_127_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_127_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_128_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_129_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_129_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_131_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_131_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_132_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_132_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_132_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_134_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_134_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_136_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_136_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_136_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_136_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_136_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_136_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_137_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_137_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_137_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_137_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_137_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_137_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_138_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_138_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_138_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_138_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_138_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_138_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_138_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_138_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_138_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_138_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_138_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_138_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_139_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_139_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_139_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_139_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_139_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_139_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_139_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_139_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_139_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_139_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_139_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_140_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_140_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_140_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_140_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_140_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_140_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_140_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_140_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_140_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_140_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_140_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_140_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_140_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_140_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_141_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_141_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_141_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_141_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_141_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_141_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_141_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_141_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_141_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_141_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_141_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_142_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_142_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_142_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_142_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_142_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_142_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_142_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_142_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_142_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_142_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_35 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_143_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_143_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_143_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_143_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_1192 ();
endmodule

