* NGSPICE file created from tiny_user_project.ext - technology: gf180mcuC

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_2 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__antenna abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__antenna I VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_1 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_4 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_64 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_64 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_1 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_1 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_1 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux4_1 I0 I1 I2 I3 S0 S1 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_8 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux2_2 I0 I1 S Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__filltie abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__filltie VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_1 D CLK Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_16 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_1 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_1 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_1 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_32 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_32 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_1 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_1 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_1 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_2 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_1 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_2 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_2 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_1 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_4 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__endcap abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__endcap VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_1 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_1 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_2 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and3_1 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_4 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_1 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_2 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_2 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor2_1 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffnq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffnq_1 D CLKN Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and4_1 A1 A2 A3 A4 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or3_1 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_1 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_2 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai222_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai222_1 A1 A2 B1 B2 C1 C2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_1 A1 A2 A3 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_2 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_1 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or4_1 A1 A2 A3 A4 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi222_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi222_1 A1 A2 B1 B2 C1 C2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__tiel abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__tiel ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_2 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai32_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai32_1 A1 A2 A3 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_20 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_20 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_4 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_2 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_12 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_12 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_2 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_4 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_2 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_2 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor3_1 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_2 A1 A2 A3 A4 ZN VDD VSS
.ends

.subckt tiny_user_project io_in[0] io_in[10] io_in[11] io_in[12] io_in[13] io_in[14]
+ io_in[15] io_in[16] io_in[17] io_in[18] io_in[19] io_in[1] io_in[20] io_in[21] io_in[22]
+ io_in[23] io_in[24] io_in[25] io_in[26] io_in[27] io_in[28] io_in[29] io_in[2] io_in[30]
+ io_in[31] io_in[32] io_in[33] io_in[34] io_in[35] io_in[36] io_in[37] io_in[3] io_in[4]
+ io_in[5] io_in[6] io_in[7] io_in[8] io_in[9] io_oeb[0] io_oeb[10] io_oeb[11] io_oeb[12]
+ io_oeb[13] io_oeb[14] io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18] io_oeb[19] io_oeb[1]
+ io_oeb[20] io_oeb[21] io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25] io_oeb[26] io_oeb[27]
+ io_oeb[28] io_oeb[29] io_oeb[2] io_oeb[30] io_oeb[31] io_oeb[32] io_oeb[33] io_oeb[34]
+ io_oeb[35] io_oeb[36] io_oeb[37] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7]
+ io_oeb[8] io_oeb[9] io_out[0] io_out[10] io_out[11] io_out[12] io_out[13] io_out[14]
+ io_out[15] io_out[16] io_out[17] io_out[18] io_out[19] io_out[1] io_out[20] io_out[21]
+ io_out[22] io_out[23] io_out[24] io_out[25] io_out[26] io_out[27] io_out[28] io_out[29]
+ io_out[2] io_out[30] io_out[31] io_out[32] io_out[33] io_out[34] io_out[35] io_out[36]
+ io_out[37] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7] io_out[8] io_out[9]
+ la_data_in[0] la_data_in[10] la_data_in[11] la_data_in[12] la_data_in[13] la_data_in[14]
+ la_data_in[15] la_data_in[16] la_data_in[17] la_data_in[18] la_data_in[19] la_data_in[1]
+ la_data_in[20] la_data_in[21] la_data_in[22] la_data_in[23] la_data_in[24] la_data_in[25]
+ la_data_in[26] la_data_in[27] la_data_in[28] la_data_in[29] la_data_in[2] la_data_in[30]
+ la_data_in[31] la_data_in[32] la_data_in[33] la_data_in[34] la_data_in[35] la_data_in[36]
+ la_data_in[37] la_data_in[38] la_data_in[39] la_data_in[3] la_data_in[40] la_data_in[41]
+ la_data_in[42] la_data_in[43] la_data_in[44] la_data_in[45] la_data_in[46] la_data_in[47]
+ la_data_in[48] la_data_in[49] la_data_in[4] la_data_in[50] la_data_in[51] la_data_in[52]
+ la_data_in[53] la_data_in[54] la_data_in[55] la_data_in[56] la_data_in[57] la_data_in[58]
+ la_data_in[59] la_data_in[5] la_data_in[60] la_data_in[61] la_data_in[62] la_data_in[63]
+ la_data_in[6] la_data_in[7] la_data_in[8] la_data_in[9] la_data_out[0] la_data_out[10]
+ la_data_out[11] la_data_out[12] la_data_out[13] la_data_out[14] la_data_out[15]
+ la_data_out[16] la_data_out[17] la_data_out[18] la_data_out[19] la_data_out[1] la_data_out[20]
+ la_data_out[21] la_data_out[22] la_data_out[23] la_data_out[24] la_data_out[25]
+ la_data_out[26] la_data_out[27] la_data_out[28] la_data_out[29] la_data_out[2] la_data_out[30]
+ la_data_out[31] la_data_out[32] la_data_out[33] la_data_out[34] la_data_out[35]
+ la_data_out[36] la_data_out[37] la_data_out[38] la_data_out[39] la_data_out[3] la_data_out[40]
+ la_data_out[41] la_data_out[42] la_data_out[43] la_data_out[44] la_data_out[45]
+ la_data_out[46] la_data_out[47] la_data_out[48] la_data_out[49] la_data_out[4] la_data_out[50]
+ la_data_out[51] la_data_out[52] la_data_out[53] la_data_out[54] la_data_out[55]
+ la_data_out[56] la_data_out[57] la_data_out[58] la_data_out[59] la_data_out[5] la_data_out[60]
+ la_data_out[61] la_data_out[62] la_data_out[63] la_data_out[6] la_data_out[7] la_data_out[8]
+ la_data_out[9] la_oenb[0] la_oenb[10] la_oenb[11] la_oenb[12] la_oenb[13] la_oenb[14]
+ la_oenb[15] la_oenb[16] la_oenb[17] la_oenb[18] la_oenb[19] la_oenb[1] la_oenb[20]
+ la_oenb[21] la_oenb[22] la_oenb[23] la_oenb[24] la_oenb[25] la_oenb[26] la_oenb[27]
+ la_oenb[28] la_oenb[29] la_oenb[2] la_oenb[30] la_oenb[31] la_oenb[32] la_oenb[33]
+ la_oenb[34] la_oenb[35] la_oenb[36] la_oenb[37] la_oenb[38] la_oenb[39] la_oenb[3]
+ la_oenb[40] la_oenb[41] la_oenb[42] la_oenb[43] la_oenb[44] la_oenb[45] la_oenb[46]
+ la_oenb[47] la_oenb[48] la_oenb[49] la_oenb[4] la_oenb[50] la_oenb[51] la_oenb[52]
+ la_oenb[53] la_oenb[54] la_oenb[55] la_oenb[56] la_oenb[57] la_oenb[58] la_oenb[59]
+ la_oenb[5] la_oenb[60] la_oenb[61] la_oenb[62] la_oenb[63] la_oenb[6] la_oenb[7]
+ la_oenb[8] la_oenb[9] user_clock2 user_irq[0] user_irq[1] user_irq[2] vdd vss wb_clk_i
+ wb_rst_i wbs_ack_o wbs_adr_i[0] wbs_adr_i[10] wbs_adr_i[11] wbs_adr_i[12] wbs_adr_i[13]
+ wbs_adr_i[14] wbs_adr_i[15] wbs_adr_i[16] wbs_adr_i[17] wbs_adr_i[18] wbs_adr_i[19]
+ wbs_adr_i[1] wbs_adr_i[20] wbs_adr_i[21] wbs_adr_i[22] wbs_adr_i[23] wbs_adr_i[24]
+ wbs_adr_i[25] wbs_adr_i[26] wbs_adr_i[27] wbs_adr_i[28] wbs_adr_i[29] wbs_adr_i[2]
+ wbs_adr_i[30] wbs_adr_i[31] wbs_adr_i[3] wbs_adr_i[4] wbs_adr_i[5] wbs_adr_i[6]
+ wbs_adr_i[7] wbs_adr_i[8] wbs_adr_i[9] wbs_cyc_i wbs_dat_i[0] wbs_dat_i[10] wbs_dat_i[11]
+ wbs_dat_i[12] wbs_dat_i[13] wbs_dat_i[14] wbs_dat_i[15] wbs_dat_i[16] wbs_dat_i[17]
+ wbs_dat_i[18] wbs_dat_i[19] wbs_dat_i[1] wbs_dat_i[20] wbs_dat_i[21] wbs_dat_i[22]
+ wbs_dat_i[23] wbs_dat_i[24] wbs_dat_i[25] wbs_dat_i[26] wbs_dat_i[27] wbs_dat_i[28]
+ wbs_dat_i[29] wbs_dat_i[2] wbs_dat_i[30] wbs_dat_i[31] wbs_dat_i[3] wbs_dat_i[4]
+ wbs_dat_i[5] wbs_dat_i[6] wbs_dat_i[7] wbs_dat_i[8] wbs_dat_i[9] wbs_dat_o[0] wbs_dat_o[10]
+ wbs_dat_o[11] wbs_dat_o[12] wbs_dat_o[13] wbs_dat_o[14] wbs_dat_o[15] wbs_dat_o[16]
+ wbs_dat_o[17] wbs_dat_o[18] wbs_dat_o[19] wbs_dat_o[1] wbs_dat_o[20] wbs_dat_o[21]
+ wbs_dat_o[22] wbs_dat_o[23] wbs_dat_o[24] wbs_dat_o[25] wbs_dat_o[26] wbs_dat_o[27]
+ wbs_dat_o[28] wbs_dat_o[29] wbs_dat_o[2] wbs_dat_o[30] wbs_dat_o[31] wbs_dat_o[3]
+ wbs_dat_o[4] wbs_dat_o[5] wbs_dat_o[6] wbs_dat_o[7] wbs_dat_o[8] wbs_dat_o[9] wbs_sel_i[0]
+ wbs_sel_i[1] wbs_sel_i[2] wbs_sel_i[3] wbs_stb_i wbs_we_i
XFILLER_140_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12902__I0 _06086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_228_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09523__A2 _03715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09671_ _03868_ _00106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_132_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08622_ _02053_ _02928_ _02929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__14966__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13607__A1 _03309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_199_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08553_ _01949_ _02859_ _02860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09287__A1 _03528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11633__I _05229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12130__I1 mod.u_cpu.rf_ram.memory\[208\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07504_ _01787_ _01812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_211_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08484_ _02041_ mod.u_cpu.rf_ram.memory\[356\]\[1\] _02790_ _02791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_51_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_196_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12830__A2 _05721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07435_ _01560_ _01743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_126_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_250_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_195_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_211_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07366_ mod.u_cpu.rf_ram.memory\[388\]\[0\] mod.u_cpu.rf_ram.memory\[389\]\[0\] mod.u_cpu.rf_ram.memory\[390\]\[0\]
+ mod.u_cpu.rf_ram.memory\[391\]\[0\] _01673_ _01666_ _01674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_195_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09105_ net2 _03405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_175_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07297_ _01604_ _01605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__14346__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09036_ mod.u_cpu.cpu.genblk3.csr.mcause3_0\[0\] _03259_ _03340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_136_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08014__A2 _02312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14496__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13146__I0 mod.u_arbiter.i_wb_cpu_rdt\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09938_ _04067_ _04068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_89_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_252_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13846__A1 _06437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_259_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09869_ _04001_ mod.u_cpu.rf_ram.memory\[538\]\[0\] _04020_ _04021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_85_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11900_ _05415_ _00788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_133_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__14120__S _07044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12880_ _06076_ _01107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_133_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_260_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_218_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11831_ _05365_ _00769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_165_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14550_ _00404_ net3 mod.u_cpu.rf_ram.memory\[412\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_92_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11762_ _05318_ _00747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_42_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10132__I0 _04193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_242_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_202_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_199_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13501_ _06559_ _01245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_201_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10713_ _04172_ _04570_ _04603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__15121__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14023__A1 mod.u_arbiter.i_wb_cpu_rdt\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14481_ _00335_ net3 mod.u_cpu.rf_ram.memory\[447\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11693_ _05271_ mod.u_cpu.rf_ram.memory\[251\]\[1\] _05269_ _05272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_1899 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_158_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13432_ _03508_ _06511_ _06514_ _03507_ _06517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_10644_ _04556_ _00391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_6_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10435__I1 _04383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13363_ _06458_ _06459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_139_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10575_ _04498_ mod.u_cpu.rf_ram.memory\[430\]\[1\] _04508_ _04510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08073__B _02379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15271__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15102_ _00956_ net3 mod.u_cpu.rf_ram.memory\[489\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10060__A2 _04143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12314_ _03696_ _05694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_181_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13294_ _06281_ _06284_ _06391_ _06392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_142_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14839__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_170_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_1281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_15033_ _00887_ net3 mod.u_cpu.rf_ram.memory\[201\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_114_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12245_ _05635_ mod.u_cpu.rf_ram.memory\[196\]\[1\] _05646_ _05648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_177_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10199__I0 _04249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09683__I _03739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12176_ _05600_ _00879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_174_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10899__A1 _04163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13137__I0 mod.u_arbiter.i_wb_cpu_rdt\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11127_ _04847_ _04887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08299__I _01533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14989__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11058_ _03984_ _04838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_249_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_95_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_5171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_77_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_92_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10009_ _04115_ mod.u_cpu.rf_ram.memory\[516\]\[1\] _04113_ _04116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_114_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_252_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_265_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10371__I0 _04363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14817_ _00671_ net3 mod.u_cpu.rf_ram.memory\[27\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_52_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11453__I _05107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14748_ _00602_ net3 mod.u_cpu.rf_ram.memory\[313\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_60_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_71_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_232_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11871__I0 _05383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_177_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14679_ _00533_ net3 mod.u_cpu.rf_ram.memory\[348\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_162_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14369__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07220_ _01527_ _01528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_193_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__15614__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_220_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11379__A2 _05058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07151_ _01439_ _01460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__09441__A1 _03670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07378__I _01527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_195_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12328__A1 _05283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08627__S0 _02048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_259_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09744__A2 _03893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13128__I0 mod.u_arbiter.i_wb_cpu_rdt\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10532__I _04429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13828__A1 _06283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07984_ _02124_ _02282_ _02290_ _02291_ _02292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_68_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09723_ _03711_ _03788_ _03909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_86_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07507__A1 _01739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_228_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09654_ _03854_ _00103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_132_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_242_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08605_ _01738_ _02874_ _02911_ _02912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_43_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15144__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09585_ _03763_ _03800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08536_ _02730_ _02842_ _02207_ _02843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_230_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07366__S0 _01673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_196_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08467_ _02303_ mod.u_cpu.rf_ram.memory\[374\]\[1\] _02773_ _01867_ _02774_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_50_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__15294__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_211_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07418_ _01605_ _01725_ _01726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_137_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08398_ _02500_ mod.u_cpu.rf_ram.memory\[436\]\[1\] _02704_ _02705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_211_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13603__I1 _06221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11614__I0 _05208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_177_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07349_ _01532_ _01657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_137_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10707__I _04574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10360_ _04364_ _00299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_136_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11739__S _05302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_174_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09019_ mod.u_arbiter.i_wb_cpu_ibus_adr\[0\] mod.u_cpu.cpu.ctrl.pc_plus_4_cy_r _03324_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_152_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10291_ _04313_ mod.u_cpu.rf_ram.memory\[476\]\[1\] _04316_ _04318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_151_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12030_ _05498_ mod.u_cpu.rf_ram.memory\[19\]\[0\] _05503_ _05504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_88_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13819__A1 _06363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_265_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_219_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09499__A1 mod.u_cpu.cpu.immdec.imm11_7\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13981_ _06946_ _06948_ _01336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_24_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3010 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_234_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12932_ _06110_ _01125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_111_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_247_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3021 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3032 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3043 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_261_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3054 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12863_ _05786_ _06064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3065 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_222_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13047__A2 _05387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3076 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_185_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08068__B _02375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3087 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3098 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14602_ _00456_ net3 mod.u_cpu.rf_ram.memory\[386\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_226_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_215_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11814_ _05354_ _00763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15582_ _01353_ net3 mod.u_arbiter.i_wb_cpu_dbus_dat\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__14511__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12794_ _06019_ mod.u_cpu.rf_ram.memory\[130\]\[1\] _06015_ _06020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__15637__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_215_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14533_ _00387_ net3 mod.u_cpu.rf_ram.memory\[421\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_109_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_214_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_11745_ _05265_ _05306_ _05307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_159_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_202_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_202_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_187_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07521__I1 mod.u_cpu.rf_ram.memory\[329\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14464_ _00318_ net3 mod.u_cpu.rf_ram.memory\[455\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11676_ _05243_ mod.u_cpu.rf_ram.memory\[256\]\[0\] _05259_ _05260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_202_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_202_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12558__A1 _05657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14661__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08515__C _02764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10408__I1 _04396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13415_ _06354_ mod.u_cpu.rf_ram.memory\[139\]\[1\] _06503_ _06505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_10627_ _04546_ _00384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_14395_ _00249_ net3 mod.u_cpu.rf_ram.memory\[490\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09423__A1 _03564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07198__I mod.u_cpu.raddr\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11230__A1 _04955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13346_ _06424_ _06443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_154_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10558_ _04498_ mod.u_cpu.rf_ram.memory\[433\]\[1\] _04494_ _04499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_115_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11649__S _05240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_192_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13277_ _06321_ _06373_ _06374_ _06375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__15017__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10489_ _04452_ _04453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_15016_ _00870_ net3 mod.u_cpu.rf_ram.memory\[207\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12228_ _05636_ _00895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12030__I0 _05498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09726__A2 _03911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07737__A1 _02040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_257_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12159_ _03727_ _04379_ _05589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_68_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10592__I0 _04514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15167__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_204_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13530__I0 _06581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_253_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08162__A1 _02449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_224_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_225_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_213_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_240_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_206_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09370_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[23\] _03610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_212_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08321_ _02592_ _02620_ _02627_ _01658_ _02628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_177_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11844__I0 _05366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_32_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_177_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11911__I _05422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09588__I _03739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08252_ _02559_ _02560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_177_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07203_ _01510_ _01511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_20_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08425__C _01678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08183_ _02321_ _02491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13210__A2 _06316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_192_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07134_ mod.u_cpu.cpu.immdec.imm24_20\[0\] _01438_ _01441_ _01442_ _01443_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__11221__A1 _04812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10024__A2 _04002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08076__S1 _02383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07728__A1 _01738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08160__C _02467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12721__A1 _05588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_247_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_210_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07967_ _02272_ mod.u_cpu.rf_ram.memory\[254\]\[0\] _02274_ _02252_ _02275_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_114_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11288__A1 _04746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09706_ _03895_ _03896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_114_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_216_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_261_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_229_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__14534__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07898_ _02202_ _02203_ _02205_ _02049_ _02206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__07571__I _01710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_243_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_228_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_216_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09637_ _03779_ _03820_ _03841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__10886__I1 mod.u_cpu.rf_ram.memory\[380\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_245_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07900__A1 _02196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09568_ _03704_ _03747_ _03748_ _03786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_130_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09102__B1 _03397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_208_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12788__A1 _03974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11835__I0 _05366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_180_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14684__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08519_ mod.u_cpu.rf_ram.memory\[341\]\[1\] _02826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__10638__I1 mod.u_cpu.rf_ram.memory\[420\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_212_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_196_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09499_ mod.u_cpu.cpu.immdec.imm11_7\[3\] mod.u_cpu.cpu.immdec.imm11_7\[4\] _03724_
+ _03725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_24_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09498__I _01441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11530_ _05161_ _00672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_23_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10263__A2 _04295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_212_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_208_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_196_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08335__C _01651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13588__I0 mod.u_arbiter.i_wb_cpu_dbus_adr\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11461_ _05113_ _00651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08208__A2 mod.u_cpu.rf_ram.memory\[566\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09405__A1 _03439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08839__S0 _02391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13200_ _06283_ _06285_ _06296_ _06306_ _06307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_183_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10412_ _04347_ _04400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_109_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14180_ _07081_ mod.u_cpu.rf_ram.memory\[8\]\[1\] _07083_ _07085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_11392_ _05046_ mod.u_cpu.rf_ram.memory\[300\]\[0\] _05067_ _05068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_139_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07967__A1 _02272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13131_ _06255_ _01179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_152_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10343_ _04302_ _04353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_174_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07746__I _01569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12012__I0 _05470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13062_ mod.u_cpu.rf_ram.memory\[69\]\[1\] _06005_ _06209_ _06211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_140_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10274_ _04305_ _00272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_79_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08070__C _02377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11268__I _04194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_239_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_191_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12013_ _05492_ _00824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_2_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_254_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08392__A1 _02188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_266_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_207_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11279__A1 _04852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13964_ _06920_ _06934_ _06935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10326__I0 _04330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_235_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_207_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_206_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09192__I0 mod.u_arbiter.i_wb_cpu_rdt\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09341__B1 _03401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12915_ _04955_ _04644_ _06099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_207_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14217__A1 _04025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13895_ _06581_ mod.u_cpu.rf_ram.memory\[112\]\[1\] _06882_ _06884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_62_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_222_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15634_ _01405_ net3 mod.u_cpu.cpu.state.o_cnt_r\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12846_ _03743_ _06052_ _01097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_2150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_146_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_221_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15565_ _01336_ net3 mod.u_arbiter.i_wb_cpu_dbus_dat\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_14_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_12777_ _05992_ mod.u_cpu.rf_ram.memory\[132\]\[0\] _06007_ _06008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_199_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14516_ _00370_ net3 mod.u_cpu.rf_ram.memory\[42\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11728_ _05295_ _00736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_159_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15496_ _01267_ net3 mod.u_arbiter.i_wb_cpu_dbus_adr\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_147_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_147_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14447_ _00301_ net3 mod.u_cpu.rf_ram.memory\[464\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11659_ _04973_ _05120_ _05247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12763__S _05996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_266_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_200_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_174_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14378_ _00232_ net3 mod.u_cpu.rf_ram.memory\[498\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_196_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__14407__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12951__A1 _06126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13329_ _06425_ _06402_ _06426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10801__I1 _04661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_157_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_233_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08870_ mod.u_cpu.rf_ram.memory\[552\]\[1\] mod.u_cpu.rf_ram.memory\[553\]\[1\] mod.u_cpu.rf_ram.memory\[554\]\[1\]
+ mod.u_cpu.rf_ram.memory\[555\]\[1\] _02472_ _02473_ _03177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__14557__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_229_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_215_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07821_ _02047_ _02129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_57_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15525__D _01296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10810__I _03941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07752_ mod.u_cpu.rf_ram.memory\[148\]\[0\] mod.u_cpu.rf_ram.memory\[149\]\[0\] mod.u_cpu.rf_ram.memory\[150\]\[0\]
+ mod.u_cpu.rf_ram.memory\[151\]\[0\] _02059_ _01723_ _02060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_84_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08135__A1 _02150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09183__I0 mod.u_arbiter.i_wb_cpu_rdt\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_225_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__14208__A1 _03775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07683_ _01850_ _01991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_93_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09422_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[30\] _03650_ _03655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_241_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_198_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_198_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_213_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_209_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_206_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11817__I0 _05342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09353_ _03415_ mod.u_scanchain_local.module_data_in\[56\] _03408_ mod.u_arbiter.i_wb_cpu_dbus_adr\[19\]
+ _03596_ _03597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XANTENNA__10458__S _04427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_178_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08304_ _02350_ _02611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11442__A1 _04965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09284_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[8\] mod.u_cpu.cpu.ctrl.o_ibus_adr\[5\] _03521_
+ _03532_ _03538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_166_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07110__A2 mod.u_cpu.cpu.csr_imm vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_178_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08235_ _01855_ _02543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_176_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_197_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_193_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13195__A1 _06126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08166_ mod.u_cpu.rf_ram.memory\[552\]\[0\] mod.u_cpu.rf_ram.memory\[553\]\[0\] mod.u_cpu.rf_ram.memory\[554\]\[0\]
+ mod.u_cpu.rf_ram.memory\[555\]\[0\] _02472_ _02473_ _02474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_101_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_134_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11745__A2 _05306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12942__A1 _03500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15332__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_238_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07117_ mod.u_cpu.cpu.decode.op26 _01426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_08097_ _02154_ _02405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_107_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_251_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08374__A1 _02148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15482__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10181__A1 _04238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08999_ _03301_ _03303_ _03304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_125_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_229_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08126__A1 _02365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_91_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_249_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10961_ _04746_ _04770_ _04771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_56_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08677__A2 mod.u_cpu.rf_ram.memory\[214\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__13670__A2 _06657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_204_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12700_ _05938_ mod.u_cpu.rf_ram.memory\[140\]\[1\] _05956_ _05958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_95_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_204_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_204_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13680_ _06689_ _06690_ _06691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_70_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10892_ _04724_ _00471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_44_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_203_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11808__I0 _05350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12631_ _05870_ _03886_ _05912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_58_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__12647__I _05873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_245_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08429__A2 mod.u_cpu.rf_ram.memory\[404\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_197_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13422__A2 _03668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_180_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10236__A2 _04263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15350_ _01125_ net3 mod.u_cpu.rf_ram.memory\[369\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12562_ _05865_ _01000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_223_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_197_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_223_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14301_ _00155_ net3 mod.u_cpu.rf_ram.memory\[537\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_129_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11513_ _05144_ mod.u_cpu.rf_ram.memory\[281\]\[0\] _05150_ _05151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_184_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15281_ _00039_ net4 mod.u_scanchain_local.module_data_in\[38\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_157_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_12493_ _05821_ _00975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_156_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_14232_ _00086_ net3 mod.u_cpu.rf_ram.memory\[571\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11444_ _05101_ _00646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11036__I1 mod.u_cpu.rf_ram.memory\[356\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_256_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_171_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08288__S1 _02594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13478__I _06537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12933__A1 _06062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14163_ _06062_ _06568_ _07073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11375_ _01968_ _05055_ _05056_ _00622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_164_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08601__A2 _02904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09892__S _04034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13114_ _06244_ _01173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_10326_ _04330_ mod.u_cpu.rf_ram.memory\[470\]\[1\] _04339_ _04341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_14094_ _07029_ _01368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_124_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13045_ _06199_ mod.u_cpu.rf_ram.memory\[107\]\[1\] _06197_ _06200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_152_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10257_ _04292_ _00268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_3_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_191_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07168__A2 _01459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_230_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10188_ _04217_ mod.u_cpu.rf_ram.memory\[490\]\[0\] _04243_ _04244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_39_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_266_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_254_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14996_ _00850_ net3 mod.u_cpu.rf_ram.memory\[65\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_93_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_207_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13110__A1 _03960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13947_ _03430_ _03433_ _06921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__08668__A2 mod.u_cpu.rf_ram.memory\[216\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_235_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13661__A2 _06404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_223_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_228_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15205__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13878_ _06422_ _06864_ _06866_ _06811_ _06870_ _01311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_50_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_250_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15617_ _01388_ net3 mod.u_cpu.rf_ram.memory\[90\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12829_ _06042_ _01090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_34_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__12472__I0 _05807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15548_ _01319_ net3 mod.u_cpu.cpu.bne_or_bge vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_188_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_187_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15355__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10077__I _04025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15479_ _01251_ net3 mod.u_cpu.rf_ram.memory\[129\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08691__I2 mod.u_cpu.rf_ram.memory\[202\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_198_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08020_ _02297_ mod.u_cpu.rf_ram.memory\[116\]\[0\] _02327_ _02328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_129_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_239_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09971_ _03762_ _04090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07319__C _01582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_258_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08922_ _02527_ mod.u_cpu.rf_ram.memory\[540\]\[1\] _03228_ _03229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10538__I0 _04481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07159__A2 mod.u_cpu.cpu.immdec.imm19_12_20\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08356__A1 _02631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_170_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08853_ _01608_ mod.u_cpu.rf_ram.memory\[38\]\[1\] _03159_ _02212_ _03160_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_131_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10163__A1 _04223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_257_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_242_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_69_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07804_ mod.u_cpu.rf_ram.memory\[173\]\[0\] _02112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_3609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08784_ mod.u_cpu.rf_ram.memory\[84\]\[1\] mod.u_cpu.rf_ram.memory\[85\]\[1\] mod.u_cpu.rf_ram.memory\[86\]\[1\]
+ mod.u_cpu.rf_ram.memory\[87\]\[1\] _01857_ _02054_ _03091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__08108__A1 _02405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09305__B1 _03555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_226_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2908 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07735_ _02042_ _02043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_2919 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_226_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07666_ _01956_ _01959_ _01973_ _01812_ _01974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__08945__I _01440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_198_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09405_ _03439_ mod.u_scanchain_local.module_data_in\[64\] _03641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_129_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_240_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07597_ _01875_ mod.u_cpu.rf_ram.memory\[356\]\[0\] _01904_ _01905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_41_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_179_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09336_ _03578_ _03582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_222_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_55_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_205_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_205_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09267_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[6\] _03524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_224_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08831__A2 _03134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12215__I0 _05605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14722__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11018__I1 mod.u_cpu.rf_ram.memory\[35\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08218_ _02084_ _02526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__13707__A3 _06714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09198_ _03471_ _00027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_193_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12915__A1 _04955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08149_ _01634_ _02457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_119_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_175_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07296__I _01603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12391__A2 _04142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11160_ _04896_ mod.u_cpu.rf_ram.memory\[337\]\[1\] _04907_ _04909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_106_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14872__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11747__S _05306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10111_ _04178_ mod.u_cpu.rf_ram.memory\[501\]\[1\] _04185_ _04188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_106_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11091_ _04796_ _04862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_248_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09217__S _03479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10042_ _01612_ _04138_ _04139_ _00206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_121_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_103_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_88_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_195_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13891__A2 _06881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08442__S1 _02748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14850_ _00704_ net3 mod.u_cpu.rf_ram.memory\[262\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_236_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15228__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09147__I0 mod.u_arbiter.i_wb_cpu_rdt\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14140__I0 _07057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13801_ _06789_ _06774_ _06800_ _06801_ _01303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__07570__A2 mod.u_cpu.rf_ram.memory\[372\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_263_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14781_ _00635_ net3 mod.u_cpu.rf_ram.memory\[297\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_4899 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11993_ _05470_ mod.u_cpu.rf_ram.memory\[569\]\[0\] _05478_ _05479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_91_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_205_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13732_ _06722_ _06657_ _06737_ _06738_ _01297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_147_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11654__A1 _04831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10944_ _04758_ _04759_ _04760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_72_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_204_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_232_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_232_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_205_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14252__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15378__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13663_ _06661_ _06369_ _06675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10098__S _04174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_204_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10875_ _04703_ _04713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_16_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_204_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_15402_ _01177_ net3 mod.u_cpu.rf_ram.memory\[359\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_220_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_12614_ _05283_ _05900_ _05901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08791__S _01517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13594_ mod.u_arbiter.i_wb_cpu_dbus_adr\[29\] mod.u_arbiter.i_wb_cpu_dbus_adr\[30\]
+ _06614_ _06618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XPHY_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_15333_ _01108_ net3 mod.u_cpu.rf_ram.memory\[99\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_12545_ _05854_ _00994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_185_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08822__A2 _03125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_177_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__12206__I0 _05609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15264_ _00021_ net4 mod.u_arbiter.i_wb_cpu_rdt\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12476_ _02535_ _05809_ _05810_ _00969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_32_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14215_ _03735_ mod.u_cpu.rf_ram.memory\[259\]\[1\] _07103_ _07105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_144_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11427_ _05071_ mod.u_cpu.rf_ram.memory\[294\]\[0\] _05090_ _05091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_125_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15195_ _01048_ net3 mod.u_cpu.rf_ram.memory\[13\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_153_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08586__A1 _01978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14146_ _07062_ _01387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_11358_ _05044_ _00617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_152_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_193_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13936__I _06910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10309_ _04266_ _04330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_98_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14077_ _03910_ _04996_ _07018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_234_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11289_ _01921_ _04997_ _04998_ _00594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__07934__I _01604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12134__A2 _05543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13331__A1 _06424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13028_ _06184_ mod.u_cpu.rf_ram.memory\[84\]\[1\] _06187_ _06189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_117_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_239_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_266_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_255_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10940__I0 _04756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_208_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_212_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09689__I1 mod.u_cpu.rf_ram.memory\[55\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14979_ _00833_ net3 mod.u_cpu.rf_ram.memory\[5\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_75_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07520_ _01827_ _01828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_47_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_235_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08510__A1 _02664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07451_ _01758_ _01759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_222_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07602__C _01657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__14745__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_195_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07382_ mod.u_cpu.rf_ram.memory\[396\]\[0\] mod.u_cpu.rf_ram.memory\[397\]\[0\] mod.u_cpu.rf_ram.memory\[398\]\[0\]
+ mod.u_cpu.rf_ram.memory\[399\]\[0\] _01689_ _01683_ _01690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_148_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09066__A2 _03368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_206_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09121_ _03419_ _00030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_148_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09596__I _03809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09052_ _03354_ _03355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_148_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_194_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08003_ _02105_ _02292_ _02310_ _02311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__08433__C _02730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_191_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14895__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_191_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10384__A1 _04230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11567__S _05184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09954_ _02547_ _04078_ _04079_ _00178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_103_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08329__A1 _02421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07844__I _02126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13322__A1 _03664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_252_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13322__B2 _06418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08905_ _02500_ _03211_ _03212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09885_ _04018_ mod.u_cpu.rf_ram.memory\[536\]\[1\] _04030_ _04032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10136__A1 _03866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13873__A2 mod.u_arbiter.i_wb_cpu_rdt\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10270__I _04301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08836_ mod.u_cpu.rf_ram.memory\[48\]\[1\] mod.u_cpu.rf_ram.memory\[49\]\[1\] mod.u_cpu.rf_ram.memory\[50\]\[1\]
+ mod.u_cpu.rf_ram.memory\[51\]\[1\] _02421_ _02393_ _03143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_218_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10931__I0 _04728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_211_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14275__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_245_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08767_ _02303_ _03073_ _03074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_85_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_174_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15520__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08188__S0 _02494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11636__A1 _04821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07718_ _01757_ _02026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08698_ mod.u_cpu.rf_ram.memory\[199\]\[1\] _03005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__13514__C _06568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07935__S0 _02242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07649_ _01919_ _01957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_241_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13389__A1 _06377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10660_ _04560_ mod.u_cpu.rf_ram.memory\[416\]\[1\] _04565_ _04567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_90_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09057__A2 mod.u_cpu.cpu.csr_imm vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_179_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09319_ _03497_ _03568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_22_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14118__S _07044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08804__A2 mod.u_cpu.rf_ram.memory\[70\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10591_ _04520_ _00374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13022__S _06182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_182_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08624__B _01602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08360__S0 _01963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12330_ _05705_ _00928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_194_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10611__A2 _04534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08343__C _01821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12261_ _05645_ mod.u_cpu.rf_ram.memory\[193\]\[0\] _05658_ _05659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_110_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_208_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_135_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08112__S0 _02403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14000_ mod.u_arbiter.i_wb_cpu_dbus_dat\[14\] _06954_ _06962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11212_ _04943_ _00572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_134_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12192_ _05334_ _05611_ _05612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xoutput7 net7 io_out[14] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_162_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_253_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11143_ _04897_ _00549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_150_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07240__A1 _01545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15050__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12116__A2 _05471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13313__A1 _06338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_249_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_5320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11074_ _04841_ mod.u_cpu.rf_ram.memory\[351\]\[1\] _04849_ _04851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_95_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_5331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14618__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10180__I _03910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14902_ _00756_ net3 mod.u_cpu.rf_ram.memory\[233\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_88_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10025_ mod.u_cpu.rf_ram.memory\[513\]\[0\] _03925_ _04126_ _04127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_5364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_49_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_209_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08740__A1 _03017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14833_ _00687_ net3 mod.u_cpu.rf_ram.memory\[271\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_5_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3940 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3951 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3962 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14764_ _00618_ net3 mod.u_cpu.rf_ram.memory\[305\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__14768__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3973 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12675__I0 _05934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3984 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11976_ _02458_ _05466_ _05467_ _00812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_60_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3995 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_232_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_229_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13715_ mod.u_cpu.cpu.immdec.imm19_12_20\[5\] _06722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_32_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_205_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10927_ _04739_ mod.u_cpu.rf_ram.memory\[373\]\[1\] _04745_ _04748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_45_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_204_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14695_ _00549_ net3 mod.u_cpu.rf_ram.memory\[340\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_147_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_108_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_205_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13646_ _06655_ _06658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_72_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_220_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10858_ _03990_ _04700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_60_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_220_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__12835__I net5 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13577_ _06608_ _01272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_158_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10789_ _04641_ mod.u_cpu.rf_ram.memory\[395\]\[1\] _04652_ _04654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XPHY_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_157_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_200_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_15316_ mod.u_cpu.cpu.o_wdata1 net3 mod.u_cpu.rf_ram_if.wdata1_r\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10602__A2 _04225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12528_ _01574_ _05842_ _05844_ _00987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_157_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15247_ _00052_ net4 mod.u_arbiter.i_wb_cpu_rdt\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_201_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12459_ _03338_ _03668_ _03359_ _03394_ _05797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_126_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08559__A1 _01963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15178_ _01031_ net3 mod.u_cpu.rf_ram.memory\[145\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_153_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13666__I _06415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_236_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_125_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14129_ _07051_ _01381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_28_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_141_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07664__I _01686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13304__A1 _06118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12107__A2 _05553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14298__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11186__I _04905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15543__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_228_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10090__I _03821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09670_ _03847_ mod.u_cpu.rf_ram.memory\[561\]\[0\] _03867_ _03868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08731__A1 _03017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_223_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08621_ mod.u_cpu.rf_ram.memory\[140\]\[1\] mod.u_cpu.rf_ram.memory\[141\]\[1\] mod.u_cpu.rf_ram.memory\[142\]\[1\]
+ mod.u_cpu.rf_ram.memory\[143\]\[1\] _02070_ _02071_ _02928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_227_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_254_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08709__B _03015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08552_ mod.u_cpu.rf_ram.memory\[319\]\[1\] _02859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_78_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07503_ _01773_ _01805_ _01810_ _01785_ _01811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_51_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08483_ _01520_ _02789_ _02790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07837__A3 _02144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_223_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07434_ _01741_ _01742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_161_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09039__A2 _01452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_189_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_211_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07365_ _01672_ _01673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_206_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_241_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09104_ _03403_ _03404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_164_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13791__A1 _06791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07296_ _01603_ _01604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_148_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09035_ _03338_ mod.u_cpu.cpu.genblk3.csr.mcause31 _03339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__15073__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09598__I0 _03802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_163_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07222__A1 _01505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07574__I _01749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_266_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08970__A1 mod.u_cpu.cpu.bufreg2.i_cnt_done vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09937_ _04066_ _04067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_131_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_217_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_219_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13846__A2 _06662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_258_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09868_ _03797_ _04003_ _04020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14910__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09770__I0 _03936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07376__I2 mod.u_cpu.rf_ram.memory\[394\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08819_ mod.u_cpu.rf_ram.memory\[31\]\[1\] _03126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_3214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_133_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09799_ _03968_ _03969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_100_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11830_ _05364_ mod.u_cpu.rf_ram.memory\[39\]\[1\] _05362_ _05365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_2_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_199_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11761_ _05304_ mod.u_cpu.rf_ram.memory\[239\]\[1\] _05316_ _05318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_199_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_260_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_158_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_199_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13500_ _03642_ _06557_ _06558_ _03648_ _06559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_1867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10712_ _04602_ _00413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_199_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14480_ _00334_ net3 mod.u_cpu.rf_ram.memory\[447\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11692_ _05249_ _05271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_202_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_158_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13431_ _06516_ _01218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__12034__A1 _03728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10643_ mod.u_cpu.rf_ram.memory\[41\]\[1\] _04532_ _04554_ _04556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_201_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08789__A1 _01493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07749__I _01487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_210_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15416__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13362_ _06391_ _06458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_195_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10574_ _04509_ _00368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_167_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10596__A1 _04242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_177_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_154_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08073__C _02380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15101_ _00955_ net3 mod.u_cpu.rf_ram.memory\[175\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_155_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12313_ _05693_ _00923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12591__S _05883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07461__A1 _01742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13293_ mod.u_arbiter.i_wb_cpu_rdt\[9\] mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat\[9\]
+ _03499_ _06391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_182_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15032_ _00886_ net3 mod.u_cpu.rf_ram.memory\[201\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_177_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12244_ _05647_ _00900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_6_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_257_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10199__I1 mod.u_cpu.rf_ram.memory\[48\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14440__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15566__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12175_ _05583_ mod.u_cpu.rf_ram.memory\[76\]\[1\] _05598_ _05600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_29_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10899__A2 _04709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11126_ _04886_ _00543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_151_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_218_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11057_ _04837_ _00523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11848__A1 _04014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14590__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12896__I0 _06086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_231_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10008_ _04090_ _04115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_5194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_209_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_264_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_149_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_266_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_236_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_218_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14816_ _00670_ net3 mod.u_cpu.rf_ram.memory\[27\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_184_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12648__I0 _05923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_149_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_264_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_252_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_233_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08248__C _02555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_205_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14747_ _00601_ net3 mod.u_cpu.rf_ram.memory\[314\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11959_ _05442_ mod.u_cpu.rf_ram.memory\[529\]\[0\] _05456_ _05457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12766__S _06000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_178_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13470__B1 _06540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_205_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_220_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14678_ _00532_ net3 mod.u_cpu.rf_ram.memory\[348\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11871__I1 mod.u_cpu.rf_ram.memory\[72\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_189_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_149_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_13629_ _06332_ _06642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_73_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_193_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13073__I0 _06217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07659__I _01758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_186_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09816__I1 _03925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15096__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13773__A1 _06309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07150_ _01458_ _01459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_158_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12820__I0 _06035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09441__A2 _03403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_172_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_201_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12328__A2 _05703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08627__S1 _02086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_236_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07394__I _01701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14933__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07983_ _01533_ _02291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_102_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_259_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13828__A2 _06824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09722_ _03908_ _00117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_132_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_256_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08704__A1 _01486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09653_ _03832_ mod.u_cpu.rf_ram.memory\[563\]\[1\] _03852_ _03854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_68_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08604_ _01977_ _02893_ _02910_ _02911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_55_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_255_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09584_ _03799_ _00088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12639__I0 _05907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09504__I0 mod.u_cpu.rf_ram.memory\[9\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08158__C _02465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08535_ mod.u_cpu.rf_ram.memory\[296\]\[1\] mod.u_cpu.rf_ram.memory\[297\]\[1\] mod.u_cpu.rf_ram.memory\[298\]\[1\]
+ mod.u_cpu.rf_ram.memory\[299\]\[1\] _01753_ _01916_ _02842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_70_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11311__I0 _05007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_179_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_247_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_242_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11580__S _05192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_224_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14313__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15439__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07366__S1 _01666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08466_ _01864_ _02772_ _02773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_195_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_196_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07417_ mod.u_cpu.rf_ram.memory\[405\]\[0\] _01725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_196_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_259_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08397_ _02111_ _02703_ _02704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_104_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_109_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07348_ _01483_ _01590_ _01655_ _01656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_176_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_178_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14463__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15589__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_192_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07279_ _01586_ _01587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_164_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09018_ _03259_ _03322_ _03323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_191_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10290_ _04317_ _00276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_117_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_254_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_215_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10750__A1 _04360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13819__A2 _06465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_259_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13980_ mod.u_arbiter.i_wb_cpu_rdt\[7\] _06938_ _06947_ mod.u_arbiter.i_wb_cpu_dbus_dat\[7\]
+ _06948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_77_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09499__A2 mod.u_cpu.cpu.immdec.imm11_7\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3000 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12931_ _06105_ mod.u_cpu.rf_ram.memory\[369\]\[1\] _06108_ _06110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_3011 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_246_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3022 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11554__I _05106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3033 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_207_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_218_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3044 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3055 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12862_ _06062_ _06063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_234_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3066 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_160_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3077 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11813_ _05350_ mod.u_cpu.rf_ram.memory\[49\]\[1\] _05352_ _05354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08068__C _02361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3088 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14601_ _00455_ net3 mod.u_cpu.rf_ram.memory\[387\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_265_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_160_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15581_ _01352_ net3 mod.u_arbiter.i_wb_cpu_dbus_dat\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3099 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_215_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12793_ _06018_ _06019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_1631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_199_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09120__A1 _03412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_261_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_230_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14532_ _00386_ net3 mod.u_cpu.rf_ram.memory\[421\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11744_ _04983_ _03823_ _05306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_148_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14806__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07682__A1 _01979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12007__A1 _05488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14463_ _00317_ net3 mod.u_cpu.rf_ram.memory\[456\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__13055__I0 _06205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11675_ _04838_ _05120_ _05259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07700__C _02007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13755__A1 mod.u_cpu.cpu.immdec.imm19_12_20\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13414_ _06504_ _01213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12558__A2 _05757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10626_ _04523_ mod.u_cpu.rf_ram.memory\[422\]\[0\] _04545_ _04546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_155_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14394_ _00248_ net3 mod.u_cpu.rf_ram.memory\[490\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12802__I0 _06010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13345_ _06441_ _06442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_183_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10557_ _04497_ _04498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09694__I _03885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_183_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14956__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13276_ _06300_ _06374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_170_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11369__I0 _05046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_170_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10488_ _04247_ _04452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_170_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15015_ _00869_ net3 mod.u_cpu.rf_ram.memory\[75\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12227_ _05635_ mod.u_cpu.rf_ram.memory\[119\]\[1\] _05632_ _05636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_142_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_194_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_9_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08934__A1 _02550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07737__A2 _02044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09982__I0 _04096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08103__I _01778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12158_ _03712_ _05588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_151_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11109_ _04864_ mod.u_cpu.rf_ram.memory\[345\]\[0\] _04874_ _04875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_42_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_190_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12089_ _05533_ mod.u_cpu.rf_ram.memory\[65\]\[1\] _05540_ _05542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12869__I0 _06035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_238_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13530__I1 mod.u_cpu.rf_ram.memory\[129\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11541__I0 _05159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_265_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08162__A2 _02452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_237_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_225_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14336__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_253_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_220_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_224_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09111__A1 _03410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08320_ _02611_ _02623_ _02626_ _01742_ _02627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_178_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14486__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08251_ _01757_ _02559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_123_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_193_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07389__I _01633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_242_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_220_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_193_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07202_ _01509_ _01510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13746__A1 mod.u_cpu.cpu.immdec.imm19_12_20\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_197_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08182_ _02476_ _02482_ _02488_ _02489_ _02490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_146_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07133_ _01427_ _01432_ _01442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__07425__A1 _01728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08722__B _02074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14171__A1 _03804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09109__I _03385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12721__A2 _05952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09973__I0 _04091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08013__I _01719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__15111__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11780__I0 _05311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07966_ _02180_ _02273_ _02274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08948__I _01422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_263_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09705_ _03894_ _03895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_68_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11288__A2 _04997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_228_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07897_ _02204_ mod.u_cpu.rf_ram.memory\[216\]\[0\] _02205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__11532__I0 _05162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09636_ _03840_ _00099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_56_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08784__S0 _01857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_216_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15261__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14829__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09567_ _03785_ _00085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12237__A1 _05642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_231_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_230_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_243_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09102__A1 _03383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08518_ mod.u_cpu.rf_ram.memory\[336\]\[1\] mod.u_cpu.rf_ram.memory\[337\]\[1\] mod.u_cpu.rf_ram.memory\[338\]\[1\]
+ mod.u_cpu.rf_ram.memory\[339\]\[1\] _01841_ _01844_ _02825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__12788__A2 _06011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09102__B2 _03402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11835__I1 mod.u_cpu.rf_ram.memory\[228\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09498_ _01441_ _03724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_145_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08616__C _01658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13037__I0 _06186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08449_ _02337_ _02755_ _01591_ _02756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_212_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_196_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07299__I _01539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11460_ _05108_ mod.u_cpu.rf_ram.memory\[28\]\[1\] _05111_ _05113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_183_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14979__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13588__I1 mod.u_arbiter.i_wb_cpu_dbus_adr\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11599__I0 _05199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_183_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_137_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08839__S1 _01552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10411_ _04399_ _00315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_109_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11391_ _04784_ _05058_ _05067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_165_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07967__A2 mod.u_cpu.rf_ram.memory\[254\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13130_ mod.u_arbiter.i_wb_cpu_rdt\[17\] mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat\[1\]
+ _06253_ _06255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_165_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10342_ _03850_ _04352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_151_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14162__A1 _03363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13061_ _02353_ _06209_ _06210_ _01154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08216__I0 mod.u_cpu.rf_ram.memory\[512\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10273_ _04298_ mod.u_cpu.rf_ram.memory\[478\]\[0\] _04304_ _04305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_3_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_155_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12012_ _05470_ mod.u_cpu.rf_ram.memory\[57\]\[0\] _05491_ _05492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_152_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_78_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_61_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_215_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14359__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15604__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_253_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13963_ _03444_ _05794_ _06934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_247_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11523__I0 _05144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11284__I _03769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10326__I1 mod.u_cpu.rf_ram.memory\[470\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09341__A1 _03386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_219_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_207_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12914_ _06098_ _01119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_207_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13894_ _06883_ _01314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__14217__A2 _05263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_235_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15633_ _01404_ net3 mod.u_cpu.cpu.state.o_cnt_r\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12845_ _01478_ _06052_ _01096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_2151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_206_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_185_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13976__A1 mod.u_arbiter.i_wb_cpu_rdt\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_203_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15564_ _01335_ net3 mod.u_arbiter.i_wb_cpu_dbus_dat\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__13976__B2 mod.u_arbiter.i_wb_cpu_dbus_dat\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12776_ _03960_ _05978_ _06007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_159_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08526__C _01887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11727_ _05289_ mod.u_cpu.rf_ram.memory\[242\]\[0\] _05294_ _05295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_148_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14515_ _00369_ net3 mod.u_cpu.rf_ram.memory\[430\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__13028__I0 _06184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_261_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_203_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15495_ _01266_ net3 mod.u_arbiter.i_wb_cpu_dbus_adr\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_30_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_230_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_202_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11658_ _05246_ _00715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_14446_ _00300_ net3 mod.u_cpu.rf_ram.memory\[464\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_174_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10609_ _04533_ _00379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07407__A1 _01709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14377_ _00231_ net3 mod.u_cpu.rf_ram.memory\[4\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_156_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11589_ _05199_ mod.u_cpu.rf_ram.memory\[268\]\[0\] _05200_ _05201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_155_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12951__A2 _03424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13328_ _06298_ _06304_ _06425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_155_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15134__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13259_ _05787_ _06356_ _06357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_115_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10014__I0 _04117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13900__A1 _06677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_123_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10714__A1 _04542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08383__A2 _02689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07820_ mod.u_cpu.rf_ram.memory\[160\]\[0\] mod.u_cpu.rf_ram.memory\[161\]\[0\] mod.u_cpu.rf_ram.memory\[162\]\[0\]
+ mod.u_cpu.rf_ram.memory\[163\]\[0\] _02125_ _02127_ _02128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_96_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15284__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_245_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07751_ _02058_ _02059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__12467__A1 _05649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07605__C _01482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08135__A2 _02435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07682_ _01979_ _01980_ _01988_ _01989_ _01990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_37_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09421_ _03496_ mod.u_scanchain_local.module_data_in\[67\] _03654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_65_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_213_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_212_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_225_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08518__S0 _01841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09352_ _03593_ _03595_ _03488_ _03596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11817__I1 mod.u_cpu.rf_ram.memory\[230\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_209_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08303_ mod.u_cpu.rf_ram.memory\[472\]\[1\] mod.u_cpu.rf_ram.memory\[473\]\[1\] mod.u_cpu.rf_ram.memory\[474\]\[1\]
+ mod.u_cpu.rf_ram.memory\[475\]\[1\] _02593_ _02454_ _02610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_100_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07646__A1 _01918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_221_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13019__I0 _06107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09283_ _03528_ _03534_ _03537_ _00048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_178_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08234_ _01688_ _02542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_21_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08165_ _02388_ _02473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_165_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07847__I _02154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_174_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07116_ mod.u_cpu.cpu.decode.op21 _01420_ _01424_ _01425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_180_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08071__A1 _02149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12942__A2 mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08096_ mod.u_cpu.rf_ram.memory\[16\]\[0\] mod.u_cpu.rf_ram.memory\[17\]\[0\] mod.u_cpu.rf_ram.memory\[18\]\[0\]
+ mod.u_cpu.rf_ram.memory\[19\]\[0\] _02403_ _02367_ _02404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_118_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__14144__A1 _03796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_175_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_216_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14501__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15627__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09571__A1 _03786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08998_ _03276_ _03302_ _03261_ _03303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_88_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07582__I _01487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_217_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_235_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07949_ mod.u_cpu.rf_ram.memory\[240\]\[0\] mod.u_cpu.rf_ram.memory\[241\]\[0\] mod.u_cpu.rf_ram.memory\[242\]\[0\]
+ mod.u_cpu.rf_ram.memory\[243\]\[0\] _02242_ _02172_ _02257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__12458__A1 mod.u_arbiter.i_wb_cpu_dbus_dat\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14651__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_229_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08126__A2 _02426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10960_ _04369_ _04713_ _04770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_56_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_217_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09874__A2 _03786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07885__A1 _01682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09619_ _03745_ _03820_ _03827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_182_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10891_ mod.u_cpu.rf_ram.memory\[37\]\[1\] _04661_ _04722_ _04724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_231_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__15007__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_188_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_12630_ _05911_ _01022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_54_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_70_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_262_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12561_ _05858_ mod.u_cpu.rf_ram.memory\[161\]\[1\] _05863_ _05865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_238_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11512_ _04873_ _05149_ _05150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_14300_ _00154_ net3 mod.u_cpu.rf_ram.memory\[537\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_15280_ _00038_ net4 mod.u_scanchain_local.module_data_in\[37\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_180_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12492_ _05813_ mod.u_cpu.rf_ram.memory\[170\]\[0\] _05820_ _05821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__15157__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_200_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14231_ _00085_ net3 mod.u_cpu.rf_ram.memory\[572\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11443_ _05096_ mod.u_cpu.rf_ram.memory\[291\]\[0\] _05100_ _05101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_137_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12933__A2 _03669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14162_ _03363_ _06631_ _07072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_11374_ _05022_ _05055_ _05056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_109_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10944__A1 _04758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13113_ _06237_ mod.u_cpu.rf_ram.memory\[100\]\[1\] _06242_ _06244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_10325_ _04340_ _00288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_14093_ _07028_ mod.u_cpu.rf_ram.memory\[245\]\[1\] _07025_ _07029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_113_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_153_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09972__I _04090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13044_ _06104_ _06199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_124_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10256_ _04276_ mod.u_cpu.rf_ram.memory\[480\]\[0\] _04291_ _04292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_79_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__12697__A1 _03904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_266_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_266_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10187_ _04242_ _04234_ _04243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_79_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_227_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07425__C _01732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14995_ _00849_ net3 mod.u_cpu.rf_ram.memory\[212\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_59_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13110__A2 _06223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_208_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_208_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_207_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13946_ _06912_ _06920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_19_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13661__A3 _06402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_235_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07876__A1 _02174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_235_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_61_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13249__I0 _06276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12838__I _05720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13877_ mod.u_cpu.cpu.immdec.imm24_20\[3\] _06867_ _06869_ _06870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_207_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13949__A1 _03438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15616_ _01387_ net3 mod.u_cpu.rf_ram.memory\[90\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12828_ _06038_ mod.u_cpu.rf_ram.memory\[125\]\[1\] _06040_ _06042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_72_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09212__I _03414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_188_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_203_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07628__A1 _01934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15547_ _01318_ net3 mod.u_cpu.cpu.decode.co_ebreak vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12759_ _04668_ _05978_ _05996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_37_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_198_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_129_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15478_ _01250_ net3 mod.u_cpu.cpu.bufreg.lsb\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_147_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_200_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_163_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10294__S _04319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14429_ _00283_ net3 mod.u_cpu.rf_ram.memory\[473\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12573__I _05709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_198_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14524__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_200_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_155_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11983__I0 _05470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_235_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09970_ _04089_ _00184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_171_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09928__I0 _04054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08921_ _02528_ _03227_ _03228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_131_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14674__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10538__I1 mod.u_cpu.rf_ram.memory\[436\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08356__A2 _02662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08852_ _02190_ _03158_ _03159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_44_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07803_ _02047_ _02111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_258_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_217_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08783_ _02051_ _03089_ _03090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_57_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08108__A2 _02409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09305__A1 _03554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07734_ _01499_ _02042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_26_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2909 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_241_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_214_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07665_ _01961_ _01966_ _01971_ _01972_ _01973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_168_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_198_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_213_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09404_ mod.u_arbiter.i_wb_cpu_dbus_adr\[27\] _03615_ _03639_ _03640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_213_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07596_ _01759_ _01903_ _01904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_80_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_197_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13404__A3 _06497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07619__A1 _01507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09335_ _03546_ _03580_ _03581_ _00057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_200_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_181_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_194_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_244_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_21_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09266_ _03506_ _03522_ _03523_ _00045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_194_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08217_ _02454_ _02525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_193_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12215__I1 mod.u_cpu.rf_ram.memory\[198\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09197_ mod.u_arbiter.i_wb_cpu_rdt\[24\] mod.u_arbiter.i_wb_cpu_dbus_dat\[21\] _03469_
+ _03471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_147_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08148_ _02129_ _02456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12915__A2 _04644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_174_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08079_ mod.u_cpu.rf_ram.memory\[0\]\[0\] mod.u_cpu.rf_ram.memory\[1\]\[0\] mod.u_cpu.rf_ram.memory\[2\]\[0\]
+ mod.u_cpu.rf_ram.memory\[3\]\[0\] _02385_ _02386_ _02387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_84_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10110_ _01594_ _04185_ _04187_ _00226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_11090_ _04861_ _00532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12679__A1 _05312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_49_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_5513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10041_ _04044_ _04138_ _04139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_5524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_212_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_209_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_264_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_88_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08201__I _01682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07245__C _01552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_64_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_217_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_60_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_229_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13800_ mod.u_cpu.cpu.immdec.imm30_25\[2\] _06772_ _06416_ _06801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09147__I1 _03438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_217_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11992_ _03767_ _04026_ _05478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_14780_ _00634_ net3 mod.u_cpu.rf_ram.memory\[297\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_57_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12151__I0 _05583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_217_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_13731_ mod.u_cpu.cpu.immdec.imm19_12_20\[6\] _06483_ _06709_ _06738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_10943_ _04708_ _04759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_17_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_232_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_189_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12851__A1 _06052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_189_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_147_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_182_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13662_ _06434_ _06644_ _06673_ _06674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_10874_ _04712_ _00465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_15401_ _01176_ net3 mod.u_cpu.rf_ram.memory\[359\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12613_ _05373_ _05900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_13593_ _06617_ _01279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_262_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_213_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_223_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_197_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__14547__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09967__I _03995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12544_ _05837_ mod.u_cpu.rf_ram.memory\[164\]\[1\] _05852_ _05854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_15332_ _00007_ net3 mod.u_cpu.rf_ram.regzero vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_129_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_200_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_185_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08283__A1 _02561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_200_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_184_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_8_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_200_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13489__I _06539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08804__C _02109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_185_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15263_ _00020_ net4 mod.u_arbiter.i_wb_cpu_rdt\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12475_ _05759_ _05809_ _05810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_177_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_177_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10217__I0 _04249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14214_ _07104_ _01414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_11426_ _04812_ _05089_ _05090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_172_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08035__A1 _01662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15194_ _01047_ net3 mod.u_cpu.rf_ram.memory\[13\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__14697__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14145_ _07057_ mod.u_cpu.rf_ram.memory\[90\]\[0\] _07061_ _07062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_11357_ _05032_ mod.u_cpu.rf_ram.memory\[306\]\[1\] _05042_ _05044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_158_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10308_ _04329_ _00282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_113_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_258_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_14076_ _07017_ _01362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_11288_ _04746_ _04997_ _04998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_3_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11737__I _05254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09535__A1 _03752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13027_ _06188_ _01142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13331__A2 _06370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10239_ _04267_ mod.u_cpu.rf_ram.memory\[483\]\[1\] _04278_ _04280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_67_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11342__A1 _04749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_254_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_266_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_208_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09299__B1 _03536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_187_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14978_ _00832_ net3 mod.u_cpu.rf_ram.memory\[5\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_35_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12142__I0 _05575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_223_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13929_ _06904_ mod.u_cpu.rf_ram.memory\[111\]\[1\] _06901_ _06905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_228_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12693__I1 _05622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15322__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_250_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07450_ _01757_ _01758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_35_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_223_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_211_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_241_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_204_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07381_ _01633_ _01689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__13901__B _06689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09120_ _03412_ _03415_ _03418_ _03419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__15472__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09051_ _03307_ _03354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_148_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_191_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07397__I _01704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08002_ _02293_ _02296_ _02309_ _02122_ _02310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_117_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_198_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08026__A1 _02293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_239_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11956__I0 _05450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10384__A2 _04381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09953_ _03899_ _04078_ _04079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_131_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_135_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08904_ mod.u_cpu.rf_ram.memory\[519\]\[1\] _03211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_170_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09884_ _04031_ _00156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10136__A2 _04202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11184__I1 _04819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_257_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09117__I _03279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_246_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_213_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_213_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08835_ mod.u_cpu.rf_ram.memory\[52\]\[1\] mod.u_cpu.rf_ram.memory\[53\]\[1\] mod.u_cpu.rf_ram.memory\[54\]\[1\]
+ mod.u_cpu.rf_ram.memory\[55\]\[1\] _02151_ _02152_ _03142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11583__S _05196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10931__I1 mod.u_cpu.rf_ram.memory\[372\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08766_ mod.u_cpu.rf_ram.memory\[127\]\[1\] _03073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_39_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07860__I _01586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08188__S1 _02495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07717_ _02022_ mod.u_cpu.rf_ram.memory\[268\]\[0\] _02024_ _02025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_2728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10199__S _04252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08697_ _02204_ mod.u_cpu.rf_ram.memory\[196\]\[1\] _03003_ _03004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_54_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_199_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07935__S1 _02172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07648_ _01914_ _01956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_54_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_202_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_198_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13389__A2 _03449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_186_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07579_ _01886_ _01887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13633__I0 mod.u_arbiter.i_wb_cpu_rdt\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_201_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09318_ _03567_ _00054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_178_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_220_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10590_ _04506_ mod.u_cpu.rf_ram.memory\[427\]\[0\] _04519_ _04520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_181_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_210_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_194_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09249_ _03502_ _03509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08360__S1 _02666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_182_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12260_ _05657_ _05650_ _05658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_147_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11211_ _04938_ mod.u_cpu.rf_ram.memory\[328\]\[0\] _04942_ _04943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08112__S1 _02152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09765__A1 _03834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12191_ _05432_ _05611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12941__I _06117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_218_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11142_ _04896_ mod.u_cpu.rf_ram.memory\[340\]\[1\] _04894_ _04897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07240__A2 mod.u_cpu.rf_ram.memory\[462\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09517__A1 _01461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13313__A2 _06363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11073_ _04850_ _00526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_150_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12372__I0 _05729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14901_ _00755_ net3 mod.u_cpu.rf_ram.memory\[234\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_209_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10024_ _04125_ _04002_ _04126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_7_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_209_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12589__S _05883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_236_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15345__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_209_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08740__A2 _03039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14832_ _00686_ net3 mod.u_cpu.rf_ram.memory\[271\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_64_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_263_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3930 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_252_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3941 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3952 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14763_ _00617_ net3 mod.u_cpu.rf_ram.memory\[306\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_205_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3963 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3974 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11975_ _05322_ _05466_ _05467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_229_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3985 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_147_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3996 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_232_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13714_ _03364_ _06657_ _06720_ _06721_ _01296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_44_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_72_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10686__I0 _04584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10926_ _01876_ _04745_ _04747_ _00482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__15495__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_232_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14694_ _00548_ net3 mod.u_cpu.rf_ram.memory\[340\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_205_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13721__B _06475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13645_ _06656_ _06657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_60_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10857_ _04699_ _00461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_108_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_220_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_158_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_220_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10438__I0 _04400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_82_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08256__A1 _02528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_185_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_169_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_13576_ mod.u_arbiter.i_wb_cpu_dbus_adr\[21\] mod.u_arbiter.i_wb_cpu_dbus_adr\[22\]
+ _06604_ _06608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_10788_ _04653_ _00438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_185_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08534__C _01833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15315_ mod.u_cpu.rf_ram_if.wdata1_r\[1\] net3 mod.u_cpu.rf_ram_if.wdata1_r\[0\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_200_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12527_ _05843_ _05842_ _05844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_157_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_258_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15246_ _00041_ net4 mod.u_arbiter.i_wb_cpu_rdt\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12458_ mod.u_arbiter.i_wb_cpu_dbus_dat\[5\] _05795_ _05796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_11409_ _05078_ _05062_ _05079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_158_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_236_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_126_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_15177_ _01030_ net3 mod.u_cpu.rf_ram.memory\[146\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12389_ _05745_ mod.u_cpu.rf_ram.memory\[177\]\[1\] _05743_ _05746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_114_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_193_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14128_ _07043_ mod.u_cpu.rf_ram.memory\[118\]\[0\] _07050_ _07051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_141_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_154_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_259_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13304__A2 _06300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14059_ mod.u_arbiter.i_wb_cpu_dbus_dat\[29\] _07000_ _07006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_98_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07881__S _02048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input3_I io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_239_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_228_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_255_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08620_ _02046_ _02926_ _02051_ _02927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08731__A2 _03030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14712__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_208_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08551_ _01962_ mod.u_cpu.rf_ram.memory\[316\]\[1\] _02857_ _02858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08709__C _02764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07502_ _01807_ mod.u_cpu.rf_ram.memory\[446\]\[0\] _01809_ _01783_ _01810_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__10677__I0 _04579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_251_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08495__A1 _02041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08482_ mod.u_cpu.rf_ram.memory\[357\]\[1\] _02789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_223_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07433_ _01630_ _01741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__14862__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_189_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_210_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07364_ _01671_ _01672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_149_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_148_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13350__C _06446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09103_ _03261_ _03403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_202_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_202_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_191_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13791__A2 _06714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14018__I _06963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07295_ _01495_ _01603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_163_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15218__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_191_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09034_ mod.u_cpu.cpu.bufreg2.i_cnt_done _03338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_175_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11929__I0 _05426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08460__B _01788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14242__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15368__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08970__A2 mod.u_cpu.cpu.immdec.imm31 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10281__I _04043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09936_ _03818_ _03883_ _04066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_132_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10109__A2 _04185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_219_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_98_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_218_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09867_ _04019_ _00151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_219_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08722__A2 _03019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_133_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08818_ _02302_ mod.u_cpu.rf_ram.memory\[28\]\[1\] _03124_ _03125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__13059__A1 _04107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14392__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_234_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09798_ _03967_ _03968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_85_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12806__A1 _05226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08749_ _02611_ _03052_ _03055_ _01680_ _03056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_61_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_183_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_214_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10668__I0 _04560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11760_ _02250_ _05316_ _05317_ _00746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_26_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08486__A1 _02672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08030__S0 _02249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_241_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_198_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09511__S _03729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10293__A1 _03791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10711_ _04593_ mod.u_cpu.rf_ram.memory\[408\]\[1\] _04600_ _04602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_144_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11691_ _05270_ _00724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_187_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_224_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13430_ _03492_ _06511_ _06514_ _03508_ _06516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_10642_ _04555_ _00390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12034__A2 _04955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08354__C _02660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_220_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_13361_ _06437_ _06447_ _06453_ _06456_ _06457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_139_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09986__A1 _04013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10456__I _04176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13782__A2 mod.u_arbiter.i_wb_cpu_rdt\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10573_ _04506_ mod.u_cpu.rf_ram.memory\[430\]\[0\] _04508_ _04509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_194_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10596__A2 _04507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15100_ _00954_ net3 mod.u_cpu.rf_ram.memory\[175\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09450__A3 _03265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12312_ _05692_ mod.u_cpu.rf_ram.memory\[185\]\[1\] _05690_ _05693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_259_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13292_ _06389_ _06390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07461__A2 _01748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_259_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15031_ _00885_ net3 mod.u_cpu.rf_ram.memory\[202\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12243_ _05645_ mod.u_cpu.rf_ram.memory\[196\]\[0\] _05646_ _05647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_177_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12174_ _05599_ _00878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08410__A1 _01709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11125_ _04880_ mod.u_cpu.rf_ram.memory\[343\]\[1\] _04884_ _04886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08961__A2 _03265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13298__A1 _06289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14735__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12345__I0 _05711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09980__I _04050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11056_ _04825_ mod.u_cpu.rf_ram.memory\[353\]\[1\] _04835_ _04837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09210__I0 mod.u_arbiter.i_wb_cpu_rdt\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11848__A2 _05374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_88_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10007_ _04114_ _00196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_5184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_49_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_67_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14098__I0 _07028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_266_1319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_4472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14815_ _00669_ net3 mod.u_cpu.rf_ram.memory\[280\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_4483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14885__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_51_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14746_ _00600_ net3 mod.u_cpu.rf_ram.memory\[314\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08477__A1 _02027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11958_ _05047_ _04118_ _05456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_17_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10909_ _04720_ mod.u_cpu.rf_ram.memory\[376\]\[1\] _04734_ _04736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_14677_ _00531_ net3 mod.u_cpu.rf_ram.memory\[34\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_149_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11889_ _05407_ _00785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_220_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11750__I _05309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13628_ _06640_ _06641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13222__A1 _06328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_242_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_192_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13559_ _06598_ _01264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_157_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_173_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_199_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_218_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_201_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14265__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15229_ _01082_ net3 mod.u_cpu.rf_ram.memory\[128\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__15510__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11536__A1 _05133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07982_ _02283_ _02286_ _02289_ _02141_ _02290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_86_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09721_ _03890_ mod.u_cpu.rf_ram.memory\[556\]\[1\] _03906_ _03908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09201__I0 mod.u_arbiter.i_wb_cpu_rdt\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08004__I1 mod.u_cpu.rf_ram.memory\[121\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11839__A2 _04223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11925__I _05432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08704__A2 _03010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_228_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09652_ _03853_ _00102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_80_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_227_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_216_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08603_ _02898_ _02900_ _02046_ _02909_ _02910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_09583_ _03740_ mod.u_cpu.rf_ram.memory\[570\]\[0\] _03798_ _03799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_83_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09504__I1 _03699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08534_ _02188_ _02837_ _02840_ _01833_ _02841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XTAP_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08468__A1 _01855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_224_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_223_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11311__I1 mod.u_cpu.rf_ram.memory\[313\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08465_ mod.u_cpu.rf_ram.memory\[375\]\[1\] _02772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_243_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_196_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_196_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15040__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07416_ mod.u_cpu.rf_ram.memory\[400\]\[0\] mod.u_cpu.rf_ram.memory\[401\]\[0\] mod.u_cpu.rf_ram.memory\[402\]\[0\]
+ mod.u_cpu.rf_ram.memory\[403\]\[0\] _01722_ _01723_ _01724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_211_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08396_ mod.u_cpu.rf_ram.memory\[437\]\[1\] _02703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_149_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_149_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_211_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14608__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07347_ _01591_ _01620_ _01654_ _01655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__09968__A1 _03919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_195_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10578__A2 _03919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07278_ _01532_ _01586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_136_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13587__I _03692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_191_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15190__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09017_ _03320_ mod.u_cpu.cpu.ctrl.i_iscomp _03321_ _03322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__08079__S0 _02385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14758__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_191_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12575__I0 _05874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_219_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10940__S _04754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_266_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13819__A3 _06668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10750__A2 _04623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09919_ _04055_ _00167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_120_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09499__A3 _03724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3001 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12930_ _06109_ _01124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_86_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_219_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3012 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_207_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3023 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3034 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3045 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_170_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12861_ _03338_ _06062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_262_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3056 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3067 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3078 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14600_ _00454_ net3 mod.u_cpu.rf_ram.memory\[387\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11812_ _05353_ _00762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3089 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_215_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15580_ _01351_ net3 mod.u_arbiter.i_wb_cpu_dbus_dat\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_27_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_199_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12792_ _06017_ _06018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14531_ _00385_ net3 mod.u_cpu.rf_ram.memory\[422\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09120__A2 _03415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11743_ _05305_ _00741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_226_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_159_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10387__S _04381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_199_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_202_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_230_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_230_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14462_ _00316_ net3 mod.u_cpu.rf_ram.memory\[456\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11674_ _05258_ _00719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07682__A2 _01980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14288__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10018__A1 _03975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10186__I _03918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13413_ _06351_ mod.u_cpu.rf_ram.memory\[139\]\[0\] _06503_ _06504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_168_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13755__A2 _06753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15533__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10625_ _04262_ _04534_ _04545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_14393_ _00247_ net3 mod.u_cpu.rf_ram.memory\[491\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_127_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10813__I0 _04663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13344_ _06121_ _06441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_10556_ _04496_ _04497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08631__A1 _01818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_182_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10914__I _04719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_185_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_13275_ _06359_ _06360_ _06373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_142_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10487_ _04451_ _00339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_154_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_154_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15014_ _00868_ net3 mod.u_cpu.rf_ram.memory\[75\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12226_ _05634_ _05635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_194_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_155_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12157_ _05587_ _00873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_68_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12318__I0 _05696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11108_ _04873_ _04869_ _04874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_78_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12088_ _05541_ _00850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_77_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_231_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11039_ _04825_ mod.u_cpu.rf_ram.memory\[356\]\[1\] _04823_ _04826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_83_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_209_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_264_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_225_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11541__I1 mod.u_cpu.rf_ram.memory\[276\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12777__S _06007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_225_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15063__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_252_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_205_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09151__S _03442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09111__A2 mod.timer_irq vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14729_ _00583_ net3 mod.u_cpu.rf_ram.memory\[323\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_221_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07122__A1 _01428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_221_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08250_ _02541_ _02557_ _01447_ _02558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_60_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_207_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_159_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07201_ _01506_ _01509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_119_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08181_ _01717_ _02489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10096__I _04176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07132_ _01439_ _01440_ _01441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_229_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14900__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07425__A2 mod.u_cpu.rf_ram.memory\[406\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14171__A2 _05397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08925__A2 mod.u_cpu.rf_ram.memory\[542\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09973__I1 mod.u_cpu.rf_ram.memory\[522\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08481__S0 _01920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_99_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12309__I0 _05679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07965_ mod.u_cpu.rf_ram.memory\[255\]\[0\] _02273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_75_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_256_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09704_ _03702_ _03883_ _03894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_74_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08689__A1 _02202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15406__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07896_ _01993_ _02204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_74_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11532__I1 mod.u_cpu.rf_ram.memory\[278\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10496__A1 _04457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_216_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09635_ _03832_ mod.u_cpu.rf_ram.memory\[565\]\[1\] _03838_ _03840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_255_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08784__S1 _02054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_244_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07900__A3 _02206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_231_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09566_ _03764_ mod.u_cpu.rf_ram.memory\[572\]\[1\] _03783_ _03785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12237__A2 _05641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_247_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_212_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10248__A1 _04285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09102__A2 _03387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11296__I0 _04999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08517_ _02778_ _02823_ _01788_ _02824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_130_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14430__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15556__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09497_ _03722_ _03723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__08185__B _01447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_212_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08448_ _02747_ _02754_ _02755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_169_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_208_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13737__A2 _06667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_183_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08379_ _02561_ _02682_ _02685_ _02080_ _02686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_23_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10410_ mod.u_cpu.rf_ram.memory\[457\]\[1\] _04383_ _04397_ _04399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__14580__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_221_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11390_ _05066_ _00627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_192_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_192_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10341_ _04351_ _00293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10420__A1 _01521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12960__A3 _06136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12548__I0 _05855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13060_ _05948_ _06209_ _06210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_124_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10272_ _04299_ _04303_ _04304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_105_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_254_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_12011_ _04294_ _04026_ _05491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_133_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_215_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_105_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_191_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08472__S0 _02751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_266_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15086__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13962_ _06932_ _06933_ _01332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_93_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_150_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_207_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_219_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12913_ _06086_ mod.u_cpu.rf_ram.memory\[399\]\[1\] _06096_ _06098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_98_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__12597__S _05889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_13893_ _06578_ mod.u_cpu.rf_ram.memory\[112\]\[0\] _06882_ _06883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_62_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_234_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15632_ _01403_ net3 mod.u_cpu.rf_ram.memory\[244\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12844_ _05788_ _05803_ _06052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13425__A1 net5 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_261_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08807__C _02664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13976__A2 _06938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15563_ _01334_ net3 mod.u_arbiter.i_wb_cpu_dbus_dat\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12775_ _06006_ _01072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_203_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11987__A1 _03834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_226_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14514_ _00368_ net3 mod.u_cpu.rf_ram.memory\[430\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11726_ _05293_ _05284_ _05294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14923__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08852__A1 _02190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15494_ _01265_ net3 mod.u_arbiter.i_wb_cpu_dbus_adr\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_230_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_203_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11039__I0 _04825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_187_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14445_ _00299_ net3 mod.u_cpu.rf_ram.memory\[465\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11657_ _05234_ mod.u_cpu.rf_ram.memory\[258\]\[1\] _05244_ _05246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_175_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12936__B1 _06113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08604__A1 _01977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10608_ mod.u_cpu.rf_ram.memory\[425\]\[1\] _04532_ _04529_ _04533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07407__A2 mod.u_cpu.rf_ram.memory\[414\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14376_ _00230_ net3 mod.u_cpu.rf_ram.memory\[4\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11588_ _04784_ _05191_ _05200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_122_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13327_ _06385_ _06424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_156_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10539_ _04485_ _00357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_183_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_155_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13258_ _03390_ _03672_ _06356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_170_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13955__I _06910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11676__S _05259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_237_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12209_ _04195_ _04125_ _05623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__11211__I0 _04938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10014__I1 mod.u_cpu.rf_ram.memory\[515\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09955__I1 _03929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13189_ _06282_ _06289_ _06295_ _06285_ _06296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__14303__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15429__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07591__A1 _01879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_238_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_56_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07750_ _01603_ _02058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_96_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13664__A1 _06672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12467__A2 _04437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13664__B2 _06472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_265_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07681_ _01886_ _01989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_38_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14453__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_237_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_226_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__15579__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09420_ _03623_ _03652_ _03653_ _00071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_52_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12300__S _05683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_253_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12219__A2 _04226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08518__S1 _01844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09351_ _03590_ _03594_ _03595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__09096__A1 mod.u_cpu.cpu.state.init_done vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_178_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_244_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_205_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08302_ _02040_ _02609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_21_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09282_ _03535_ mod.u_scanchain_local.module_data_in\[45\] _03536_ mod.u_arbiter.i_wb_cpu_dbus_adr\[8\]
+ _03537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__08843__A1 _02191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08233_ _02523_ _02524_ _02540_ _02469_ _02541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_220_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08164_ _02329_ _02472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_147_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09643__I0 _03832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07115_ _01423_ _01424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_146_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14026__I _06970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08095_ _01856_ _02403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_161_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14144__A2 _05397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_255_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11202__I0 _04936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09571__A2 _03788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08997_ mod.u_cpu.rf_ram_if.rdata1 _03248_ mod.u_cpu.rf_ram_if.rtrig1 _03302_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_125_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_214_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_75_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07948_ _01740_ _02241_ _02255_ _02256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_25_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13655__A1 _06304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_228_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07879_ _02149_ _02169_ _02186_ _02187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_55_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07334__A1 _01607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_216_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09618_ _03826_ _00095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08694__I _01560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13407__A1 _03790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_216_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10890_ _02427_ _04722_ _04723_ _00470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__14946__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_243_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_225_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09549_ _03770_ _03771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_197_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11969__A1 _05448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_240_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08834__A1 _01693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12560_ _05864_ _00999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_93_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_212_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_200_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11511_ _05124_ _05149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_133_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_196_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12491_ _05334_ _05767_ _05820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_138_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_200_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14230_ _00084_ net3 mod.u_cpu.rf_ram.memory\[572\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_184_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11442_ _04965_ _05089_ _05100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11373_ _04369_ _05020_ _05055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_165_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14161_ _07067_ mod.u_cpu.cpu.ctrl.i_jump _07071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_109_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08693__S0 _01578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_192_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14326__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10944__A2 _04759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13112_ _06243_ _01172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_10324_ _04326_ mod.u_cpu.rf_ram.memory\[470\]\[0\] _04339_ _04340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_3_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14092_ _06903_ _07028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_113_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12146__A1 _05187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13775__I _06776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10255_ _04290_ _04137_ _04291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_13043_ _06198_ _01148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08445__S0 _02751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09011__A1 mod.u_cpu.cpu.bufreg.lsb\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13708__C _06365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_266_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14476__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10186_ _03918_ _04242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_121_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_152_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_232_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14994_ _00848_ net3 mod.u_cpu.rf_ram.memory\[212\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_187_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_247_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_13945_ _06918_ _06919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_47_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_219_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_208_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13876_ _06868_ _06837_ _06869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_235_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15615_ _01386_ net3 mod.u_cpu.rf_ram.memory\[289\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_216_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12827_ _02313_ _06040_ _06041_ _01089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_61_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15546_ _01317_ net3 mod.u_cpu.cpu.decode.op21 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12758_ _05995_ _01066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_203_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_231_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_203_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_188_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15101__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11709_ _05271_ mod.u_cpu.rf_ram.memory\[253\]\[1\] _05280_ _05282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_203_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_202_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15477_ _01249_ net3 mod.u_cpu.cpu.bufreg.lsb\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12689_ mod.u_cpu.rf_ram.memory\[77\]\[1\] _05950_ _05947_ _05951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_175_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14428_ _00282_ net3 mod.u_cpu.rf_ram.memory\[473\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_163_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_200_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12385__A1 _05742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08272__C _02555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14359_ _00213_ net3 mod.u_cpu.rf_ram.memory\[508\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_200_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15251__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_196_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_226_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_196_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__14819__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13185__I0 mod.u_arbiter.i_wb_cpu_rdt\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08920_ mod.u_cpu.rf_ram.memory\[541\]\[1\] _03227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_130_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09928__I1 mod.u_cpu.rf_ram.memory\[52\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08436__S0 _01994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07683__I _01850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13885__A1 _06735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08851_ mod.u_cpu.rf_ram.memory\[39\]\[1\] _03158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_97_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07802_ _02109_ _02110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_111_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__13637__A1 mod.u_cpu.cpu.immdec.imm31 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08782_ mod.u_cpu.rf_ram.memory\[80\]\[1\] mod.u_cpu.rf_ram.memory\[81\]\[1\] mod.u_cpu.rf_ram.memory\[82\]\[1\]
+ mod.u_cpu.rf_ram.memory\[83\]\[1\] _02249_ _02107_ _03089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__14969__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09604__S _03815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11499__I0 _05114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07733_ _01743_ _02041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_37_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_226_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07664_ _01686_ _01972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_129_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12860__A2 mod.u_cpu.rf_ram_if.rtrig1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_92_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09403_ _03614_ _03636_ _03638_ _03639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_225_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07595_ mod.u_cpu.rf_ram.memory\[357\]\[0\] _01903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_222_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09334_ _03554_ mod.u_scanchain_local.module_data_in\[53\] _03555_ mod.u_arbiter.i_wb_cpu_dbus_adr\[16\]
+ _03581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_179_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_139_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_221_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11671__I0 _05243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09265_ _03516_ mod.u_scanchain_local.module_data_in\[42\] _03518_ mod.u_arbiter.i_wb_cpu_dbus_adr\[5\]
+ _03523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_178_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14349__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07858__I _01765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08216_ mod.u_cpu.rf_ram.memory\[512\]\[0\] mod.u_cpu.rf_ram.memory\[513\]\[0\] mod.u_cpu.rf_ram.memory\[514\]\[0\]
+ mod.u_cpu.rf_ram.memory\[515\]\[0\] _02494_ _02495_ _02524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_09196_ _03470_ _00026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_119_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_194_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08182__C _02489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11423__I0 _05087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10226__I1 _04111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08147_ _02454_ _02455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_147_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14117__A2 _03911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08078_ _01581_ _02386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_175_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14499__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10040_ _03991_ _04137_ _04138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_5514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_49_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_251_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_130_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_248_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_229_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11991_ _05477_ _00817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_112_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13730_ _06456_ _06725_ _06728_ _06736_ _06640_ _06737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_10942_ _03857_ _04758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_16_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09313__I _03413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_232_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_205_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_231_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15124__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_250_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_188_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13661_ _06309_ _06404_ _06402_ _06673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_43_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14053__A1 mod.u_arbiter.i_wb_cpu_rdt\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10873_ _04698_ mod.u_cpu.rf_ram.memory\[382\]\[1\] _04710_ _04712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_15400_ _01175_ net3 mod.u_cpu.rf_ram.memory\[0\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_12612_ _05899_ _01016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__09855__I0 _04001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13592_ mod.u_arbiter.i_wb_cpu_dbus_adr\[28\] mod.u_arbiter.i_wb_cpu_dbus_adr\[29\]
+ _06614_ _06617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_197_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_197_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15331_ _01107_ net3 mod.u_cpu.rf_ram.memory\[246\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_12543_ _05853_ _00993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09480__A1 _01461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08283__A2 _02586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__15274__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_200_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_15262_ _00018_ net4 mod.u_arbiter.i_wb_cpu_rdt\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_138_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12474_ _05395_ _04033_ _05809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08092__C _02359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14213_ _03699_ mod.u_cpu.rf_ram.memory\[259\]\[0\] _07103_ _07104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_138_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11425_ _04995_ _05089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10194__I _04247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_184_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15193_ _01046_ net3 mod.u_cpu.rf_ram.memory\[140\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08035__A2 _02342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14144_ _03796_ _05397_ _07061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11356_ _05043_ _00616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_153_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10307_ _04326_ mod.u_cpu.rf_ram.memory\[473\]\[0\] _04328_ _04329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_98_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07717__B _02024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_193_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_180_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14075_ _06904_ mod.u_cpu.rf_ram.memory\[114\]\[1\] _07015_ _07017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_11287_ _04994_ _04996_ _04997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13867__A1 _06823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11717__I1 mod.u_cpu.rf_ram.memory\[248\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09535__A2 _03758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13026_ _06186_ mod.u_cpu.rf_ram.memory\[84\]\[0\] _06187_ _06188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_10238_ _04279_ _00262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_117_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_266_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_266_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_39_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10169_ _04230_ _04229_ _04231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_79_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14977_ _00831_ net3 mod.u_cpu.rf_ram.memory\[19\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_130_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09299__A1 _03535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13928_ _06903_ _06904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_35_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_208_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09223__I _03406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_207_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_262_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_179_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13859_ _06664_ _06851_ _06852_ _06464_ _06853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_223_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_223_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_206_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_204_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07380_ _01687_ _01688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__15617__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_250_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_204_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_203_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_163_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_203_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15529_ _01300_ net3 mod.u_cpu.cpu.immdec.imm19_12_20\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_128_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_198_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09050_ _03250_ _03353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_15_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_176_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08001_ _02283_ _02301_ _02307_ _02308_ _02309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_191_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14641__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_191_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_237_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_190_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08730__C _01695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09952_ _03896_ _04077_ _04078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_131_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__14791__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08903_ _02527_ mod.u_cpu.rf_ram.memory\[516\]\[1\] _03209_ _03210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08302__I _02040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09883_ _04023_ mod.u_cpu.rf_ram.memory\[536\]\[0\] _04030_ _04031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_252_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08834_ _01693_ _03121_ _03140_ _02380_ _03141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_258_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08765_ _02297_ mod.u_cpu.rf_ram.memory\[124\]\[1\] _03071_ _03072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_73_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15147__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11663__I _05249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08458__B _02763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07716_ _01729_ _02023_ _02024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_260_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_254_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_226_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08696_ _03001_ _03002_ _03003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_54_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_213_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10279__I _04308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11892__I0 _05385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07647_ _01915_ _01945_ _01954_ _01768_ _01955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__12695__S _05953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15297__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_198_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07578_ _01532_ _01886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_167_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13633__I1 _03458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_181_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09317_ _03415_ mod.u_scanchain_local.module_data_in\[50\] _03562_ _03566_ _03567_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_178_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09462__A1 _03686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_210_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_194_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09248_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[2\] _03508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_193_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09179_ mod.u_arbiter.i_wb_cpu_rdt\[16\] mod.u_arbiter.i_wb_cpu_dbus_dat\[13\] _03459_
+ _03461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_166_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11210_ _04804_ _04926_ _04942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11021__A1 _04812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12190_ _05610_ _00883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09765__A2 _03942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11572__A2 _05188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11141_ _04879_ _04896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10742__I _04621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13849__A1 _06739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11072_ _04843_ mod.u_cpu.rf_ram.memory\[351\]\[0\] _04849_ _04850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_150_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08212__I _01489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09517__A2 _01778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07256__C _01525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_49_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14900_ _00754_ net3 mod.u_cpu.rf_ram.memory\[234\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10023_ _03979_ _04125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12372__I1 mod.u_cpu.rf_ram.memory\[499\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_49_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_264_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_5355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_102_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_48_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14831_ _00685_ net3 mod.u_cpu.rf_ram.memory\[272\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_4643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12669__I _05709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3920 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3931 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3942 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11088__A1 _04859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14762_ _00616_ net3 mod.u_cpu.rf_ram.memory\[306\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3953 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14514__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3964 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11974_ _03893_ _04108_ _05466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_17_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3975 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_205_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3986 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13713_ mod.u_cpu.cpu.immdec.imm19_12_20\[5\] _06704_ _06471_ _06693_ _06656_ _06721_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XANTENNA__11883__I0 _05385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3997 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10925_ _04746_ _04745_ _04747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_244_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_189_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14693_ _00547_ net3 mod.u_cpu.rf_ram.memory\[341\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_225_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07700__A1 _01992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_186_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_220_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13644_ _06655_ _06656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_147_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10856_ _04698_ mod.u_cpu.rf_ram.memory\[384\]\[1\] _04696_ _04699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_176_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12588__A1 _05443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__14664__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10438__I1 mod.u_cpu.rf_ram.memory\[452\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__10917__I _03827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_13575_ _06607_ _01271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_158_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10787_ _04637_ mod.u_cpu.rf_ram.memory\[395\]\[0\] _04652_ _04653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07498__I _01603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_15314_ mod.u_cpu.cpu.o_wen0 net3 mod.u_cpu.rf_ram_if.wen0_r vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12526_ _05487_ _05843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_201_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_200_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15245_ _00030_ net4 mod.u_arbiter.i_wb_cpu_rdt\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12457_ mod.u_arbiter.i_wb_cpu_dbus_dat\[4\] _05794_ _05795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_138_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13001__A2 _03353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11408_ _03712_ _05078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_15176_ _01029_ net3 mod.u_cpu.rf_ram.memory\[146\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_153_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12388_ _05710_ _05745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_67_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14127_ _03828_ _05631_ _07050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_67_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11339_ _05031_ _05032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_153_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_141_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14058_ _07003_ _07005_ _01356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_97_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13009_ _06176_ _01136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_67_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_234_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08811__S0 _02211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_254_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09154__S _03442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08550_ _01934_ _02856_ _02857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_242_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_236_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_208_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12815__A2 _06031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07501_ _01779_ _01808_ _01809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_63_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08481_ mod.u_cpu.rf_ram.memory\[352\]\[1\] mod.u_cpu.rf_ram.memory\[353\]\[1\] mod.u_cpu.rf_ram.memory\[354\]\[1\]
+ mod.u_cpu.rf_ram.memory\[355\]\[1\] _01920_ _02666_ _02788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__08495__A2 mod.u_cpu.rf_ram.memory\[332\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_223_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07432_ _01488_ _01740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_50_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11626__I0 _05208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_195_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__10827__I _04621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07363_ _01537_ _01671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09444__A1 _03353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09102_ _03383_ _03387_ _03397_ _03402_ _00008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_149_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07294_ _01492_ _01602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_175_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09033_ _03258_ _03337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_191_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_191_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12051__I0 _05498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_176_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09935_ _04065_ _00173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_113_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12503__A1 _05563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_252_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_246_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_213_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09866_ _04018_ mod.u_cpu.rf_ram.memory\[53\]\[1\] _04015_ _04019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14537__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_259_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10365__I0 _04363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07871__I _01646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08817_ _02369_ _03123_ _03124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_86_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13059__A2 _05589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09797_ _03788_ _03966_ _03967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_3216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07930__A1 _01819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10117__I0 _04178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08748_ _02585_ _03053_ _03054_ _01751_ _03055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__10003__S _04109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__12806__A2 _05320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_261_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_214_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_199_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10817__A1 _04262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_226_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__14687__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08679_ mod.u_cpu.rf_ram.memory\[210\]\[1\] mod.u_cpu.rf_ram.memory\[211\]\[1\] _01807_
+ _02986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_1825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08030__S1 _02098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09798__I _03967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10710_ _04601_ _00412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_53_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11690_ _05268_ mod.u_cpu.rf_ram.memory\[251\]\[0\] _05269_ _05270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_1869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_201_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_186_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_263_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10641_ mod.u_cpu.rf_ram.memory\[41\]\[0\] _04396_ _04554_ _04555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_195_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13360_ _06455_ _06456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_158_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_194_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08207__I _02306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09986__A2 _03851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10572_ _04218_ _04507_ _04508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_194_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07997__A1 _02303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11769__S _05321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12311_ _05634_ _05692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12990__A1 _05780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_194_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12952__I _06128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_213_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13291_ _06384_ _06385_ _06387_ _06388_ _06389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_177_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15030_ _00884_ net3 mod.u_cpu.rf_ram.memory\[202\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12242_ _05367_ _05611_ _05646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12042__I0 _05501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_181_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15312__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_194_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12173_ _05575_ mod.u_cpu.rf_ram.memory\[76\]\[0\] _05598_ _05599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_181_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11124_ _04885_ _00542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_231_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13298__A2 _06390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11055_ _04836_ _00522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_7_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_265_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10356__I0 _04348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_77_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15462__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_236_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_237_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10006_ _04096_ mod.u_cpu.rf_ram.memory\[516\]\[0\] _04113_ _04114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_5174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_225_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07921__A1 _02120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_252_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_14814_ _00668_ net3 mod.u_cpu.rf_ram.memory\[280\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_4473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_218_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_224_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_229_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_251_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14745_ _00599_ net3 mod.u_cpu.rf_ram.memory\[315\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11957_ _05455_ _00805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_44_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08477__A2 _02783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07730__B _02037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10908_ _04735_ _00476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_14676_ _00530_ net3 mod.u_cpu.rf_ram.memory\[34\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11888_ _05406_ mod.u_cpu.rf_ram.memory\[227\]\[1\] _05402_ _05407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_60_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_264_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_220_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13627_ _06415_ _06640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_38_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10839_ _04569_ _04687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_186_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_157_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13558_ mod.u_arbiter.i_wb_cpu_dbus_adr\[13\] mod.u_arbiter.i_wb_cpu_dbus_adr\[14\]
+ _06594_ _06598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12281__I0 _05662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_203_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_203_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07532__S0 _01826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12509_ _05343_ _05831_ _05832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_195_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12862__I _06062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13489_ _06539_ _06552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_201_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_15228_ _01081_ net3 mod.u_cpu.rf_ram.memory\[128\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_12_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_236_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_172_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15159_ _01012_ net3 mod.u_cpu.rf_ram.memory\[155\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08401__A2 mod.u_cpu.rf_ram.memory\[438\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_259_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07981_ _02135_ mod.u_cpu.rf_ram.memory\[102\]\[0\] _02288_ _02139_ _02289_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_234_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13289__A2 _03428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09720_ _03907_ _00116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_101_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_228_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07905__B _02212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10347__I0 _04345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11839__A3 _03753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08004__I2 mod.u_cpu.rf_ram.memory\[122\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_255_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_210_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09362__B1 _03517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09651_ _03847_ mod.u_cpu.rf_ram.memory\[563\]\[0\] _03852_ _03853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_94_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_110_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08602_ _01852_ _02901_ _02908_ _01887_ _02909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_209_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09582_ _03758_ _03797_ _03798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_83_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_243_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08533_ _02225_ _02838_ _02839_ _01683_ _02840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_70_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_208_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_70_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11472__A1 _05022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_208_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13361__C _06456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08464_ _02059_ mod.u_cpu.rf_ram.memory\[372\]\[1\] _02770_ _02771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_24_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07415_ _01500_ _01723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__09417__A1 _03614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08395_ mod.u_cpu.rf_ram.memory\[432\]\[1\] mod.u_cpu.rf_ram.memory\[433\]\[1\] mod.u_cpu.rf_ram.memory\[434\]\[1\]
+ mod.u_cpu.rf_ram.memory\[435\]\[1\] _02688_ _02475_ _02702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_149_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07346_ _01489_ _01629_ _01653_ _01654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_177_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07523__S0 _01826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13868__I _06365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12972__A1 _06142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15335__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07277_ _01572_ _01576_ _01583_ _01584_ _01585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__07866__I _02154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_178_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_163_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09016_ mod.u_cpu.cpu.state.o_cnt_r\[2\] mod.u_cpu.cpu.ctrl.i_iscomp _03321_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__12024__I0 _05498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_191_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_191_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08079__S1 _02386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11388__I _04531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12575__I1 mod.u_cpu.rf_ram.memory\[15\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_219_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__15485__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09918_ _04054_ mod.u_cpu.rf_ram.memory\[531\]\[1\] _04052_ _04055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_150_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10338__I0 _04348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_247_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_218_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08156__A1 _02462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09353__B1 _03408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09849_ _03771_ _03996_ _04007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_98_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_111_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3002 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3013 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_234_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_234_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3024 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_160_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3035 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12860_ _06060_ mod.u_cpu.rf_ram_if.rtrig1 _06061_ mod.u_cpu.rf_ram.regzero _01102_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_248_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_206_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3046 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3057 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3068 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11811_ _05342_ mod.u_cpu.rf_ram.memory\[49\]\[0\] _05352_ _05353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_2334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_233_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3079 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10668__S _04571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12791_ _05105_ _06017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_226_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_261_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14530_ _00384_ net3 mod.u_cpu.rf_ram.memory\[422\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11742_ _05304_ mod.u_cpu.rf_ram.memory\[240\]\[1\] _05302_ _05305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_215_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_199_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11463__A1 _04838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_226_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_187_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14461_ _00315_ net3 mod.u_cpu.rf_ram.memory\[457\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11673_ _05250_ mod.u_cpu.rf_ram.memory\[250\]\[1\] _05256_ _05258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_186_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_161_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13412_ _03910_ _06011_ _06503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_128_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10624_ _04544_ _00383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_139_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14392_ _00246_ net3 mod.u_cpu.rf_ram.memory\[491\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_167_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07514__S0 _01819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11499__S _05140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_183_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13343_ _06437_ _06418_ _06403_ _06439_ _06440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_10_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10555_ _03761_ _04496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_259_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07285__I3 mod.u_cpu.rf_ram.memory\[499\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07776__I _01671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14702__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13274_ _06371_ _06372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_136_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10486_ _04450_ mod.u_cpu.rf_ram.memory\[445\]\[1\] _04448_ _04451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_15013_ _00867_ net3 mod.u_cpu.rf_ram.memory\[74\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_170_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12715__A1 _03918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12225_ _05404_ _05634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_155_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_190_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12156_ _05583_ mod.u_cpu.rf_ram.memory\[206\]\[1\] _05585_ _05587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__13727__B _06321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14852__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12318__I1 mod.u_cpu.rf_ram.memory\[189\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11107_ _04024_ _04873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__12123__S _05564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12087_ _05539_ mod.u_cpu.rf_ram.memory\[65\]\[0\] _05540_ _05541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10329__I0 _04326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09195__I0 mod.u_arbiter.i_wb_cpu_rdt\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_237_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_204_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11038_ _04796_ _04825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_42_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09895__A1 _03829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_253_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15208__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_225_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09647__A1 _03788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12989_ mod.u_cpu.cpu.genblk3.csr.mcause3_0\[1\] _06161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_206_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14728_ _00582_ net3 mod.u_cpu.rf_ram.memory\[323\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_162_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_220_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__14232__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15358__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14659_ _00513_ net3 mod.u_cpu.rf_ram.memory\[358\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_127_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_221_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07200_ _01507_ _01508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_08180_ _02483_ mod.u_cpu.rf_ram.memory\[558\]\[0\] _02486_ _02487_ _02488_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_158_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_203_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12954__A1 _06125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_174_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07131_ _01437_ _01440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_174_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08622__A2 _02928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14382__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07686__I _01993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_173_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10568__I0 _04498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08511__S _01664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08481__S1 _02666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_229_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07964_ _01537_ _02272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_214_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08138__A1 _01475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09186__I0 mod.u_arbiter.i_wb_cpu_rdt\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09703_ _03724_ _03892_ _03893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_96_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07895_ mod.u_cpu.rf_ram.memory\[217\]\[0\] _02203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_68_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_216_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09634_ _02510_ _03838_ _03839_ _00098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_95_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_249_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_249_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_215_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09565_ _03784_ _00084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_24_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08516_ mod.u_cpu.rf_ram.memory\[344\]\[1\] mod.u_cpu.rf_ram.memory\[345\]\[1\] mod.u_cpu.rf_ram.memory\[346\]\[1\]
+ mod.u_cpu.rf_ram.memory\[347\]\[1\] _02751_ _02748_ _02823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__10248__A2 _04137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11296__I1 mod.u_cpu.rf_ram.memory\[316\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09496_ _03718_ _03721_ _03722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_58_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_169_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08310__A1 _02198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_196_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08447_ _02230_ _02750_ _02753_ _02754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__10287__I _03781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_211_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_208_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_168_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__12245__I0 _05635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14725__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_184_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13737__A3 _06669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08378_ _02560_ _02683_ _02684_ _02594_ _02685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_149_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07329_ _01568_ _01637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_139_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_256_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10340_ _04345_ mod.u_cpu.rf_ram.memory\[468\]\[1\] _04349_ _04351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_125_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_192_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14875__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_191_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10271_ _04302_ _04303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_180_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08377__A1 _02656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12010_ _05490_ _00823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_151_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_191_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08472__S1 _02748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_266_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_266_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08129__A1 _02157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_266_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09177__I0 _03458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13122__A1 _06249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_232_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_219_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08220__I _01538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13961_ mod.u_arbiter.i_wb_cpu_rdt\[3\] _06906_ _06928_ _03441_ _06933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_93_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09877__A1 _03996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11782__S _05331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_207_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_235_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_12912_ _06097_ _01118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_219_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_171_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13892_ _03872_ _06223_ _06882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_24_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_207_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10731__I0 _04598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_262_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14255__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15631_ _01402_ net3 mod.u_cpu.rf_ram.memory\[244\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12843_ _06051_ _01095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09629__A1 _03702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15500__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13425__A2 _03677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15562_ _01333_ net3 mod.u_arbiter.i_wb_cpu_dbus_dat\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_199_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12484__I0 _05807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12774_ mod.u_cpu.rf_ram.memory\[133\]\[1\] _06005_ _06003_ _06006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_187_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_202_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11987__A2 _04068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14513_ _00367_ net3 mod.u_cpu.rf_ram.memory\[431\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11725_ _03857_ _05293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_1474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10197__I _04250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_199_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15493_ _01264_ net3 mod.u_arbiter.i_wb_cpu_dbus_adr\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13189__A1 _06282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11039__I1 mod.u_cpu.rf_ram.memory\[356\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14444_ _00298_ net3 mod.u_cpu.rf_ram.memory\[465\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11656_ _05245_ _00714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_70_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08823__C _02185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12936__B2 _06063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10607_ _04531_ _04532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_122_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14375_ _00229_ net3 mod.u_cpu.rf_ram.memory\[500\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11587_ _05143_ _05199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08604__A2 _02893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13326_ _06130_ _06423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_128_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_196_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_183_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_171_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10538_ _04481_ mod.u_cpu.rf_ram.memory\[436\]\[1\] _04483_ _04485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_157_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_171_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12539__I1 _05765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13257_ _06355_ _01205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_10469_ _04043_ _04439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_170_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08368__A1 _01567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12208_ _03698_ _05622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__13361__A1 _06437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13188_ _06291_ _06293_ _06281_ _06294_ _06295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XANTENNA__10175__A1 _04233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_233_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_12139_ _05520_ _05575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_96_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15030__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09168__I0 mod.u_arbiter.i_wb_cpu_rdt\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09317__B1 _03562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09226__I _03488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07591__A2 mod.u_cpu.rf_ram.memory\[366\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09868__A1 _03797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_226_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11675__A1 _04838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07680_ _01981_ _01984_ _01987_ _01972_ _01988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__10722__I0 _04608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08540__A1 _01807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09162__S _03442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07194__I2 mod.u_cpu.rf_ram.memory\[450\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07974__S0 _02125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15180__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12587__I _05373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_252_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09350_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[19\] mod.u_cpu.cpu.ctrl.o_ibus_adr\[18\] _03594_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__14748__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09096__A2 _03391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08301_ _02590_ _02596_ _02102_ _02607_ _02608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_221_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_209_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09281_ _03517_ _03536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_178_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08232_ _02525_ _02531_ _02538_ _02539_ _02540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__12227__I0 _05635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14898__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_197_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08163_ _01688_ _02471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_105_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09643__I1 mod.u_cpu.rf_ram.memory\[564\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10789__I0 _04641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07114_ _01421_ _01422_ _01423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_08094_ _02348_ _02394_ _02401_ _02185_ _02402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_174_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10771__S _04638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_255_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10166__A1 _04225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_216_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_173_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_248_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08996_ _03261_ mod.u_cpu.cpu.bufreg.i_sh_signed _03300_ _01422_ _03301_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_125_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09159__I0 mod.u_arbiter.i_wb_cpu_rdt\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14152__I0 _07055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__14278__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08040__I _02347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07947_ _02170_ _02243_ _02254_ _02207_ _02255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_56_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_229_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15523__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_217_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11666__A1 _03665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07878_ _02170_ _02173_ _02184_ _02185_ _02186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_141_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_244_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07334__A2 mod.u_cpu.rf_ram.memory\[492\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09617_ _03800_ mod.u_cpu.rf_ram.memory\[567\]\[1\] _03824_ _03826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08908__C _02469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_204_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_204_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09548_ _03769_ _03770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_262_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_58_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_197_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09479_ mod.u_cpu.cpu.decode.op21 _01426_ _01440_ _03705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_200_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08834__A2 _03121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11510_ _05148_ _00665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_200_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_212_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_184_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12490_ _05819_ _00974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_71_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_200_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11441_ _05099_ _00645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09244__C1 _03408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_221_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14160_ _07070_ _01392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_11372_ _05054_ _00621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_164_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08215__I _02097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_180_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08693__S1 _01714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_180_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13111_ _06230_ mod.u_cpu.rf_ram.memory\[100\]\[0\] _06242_ _06243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_124_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10323_ _04180_ _04327_ _04339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_14091_ _02258_ _07025_ _07027_ _01367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_125_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15053__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12146__A2 _05552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13343__A1 _06437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_13042_ _06186_ mod.u_cpu.rf_ram.memory\[107\]\[0\] _06197_ _06198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_10254_ _03985_ _04290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_152_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09011__A2 _03292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08445__S1 _02748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_182_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10185_ _04241_ _00247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_67_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10952__I0 _04756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07573__A2 _01880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08770__A1 _02293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14993_ _00847_ net3 mod.u_cpu.rf_ram.memory\[64\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_208_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13944_ _06913_ _06918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_75_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10704__I0 _04593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_234_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13875_ mod.u_cpu.cpu.immdec.imm24_20\[4\] _06868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_75_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15614_ _01385_ net3 mod.u_cpu.rf_ram.memory\[289\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11409__A1 _05078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12200__I _05229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12826_ _06032_ _06040_ _06041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_62_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_250_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_203_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12757_ _05984_ mod.u_cpu.rf_ram.memory\[80\]\[1\] _05993_ _05995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_15545_ _01316_ net3 mod.u_cpu.cpu.decode.op22 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_230_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11708_ _02269_ _05280_ _05281_ _00730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_163_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10632__A2 _04548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15476_ _00006_ net3 mod.u_cpu.cpu.ctrl.pc_plus_offset_cy_r vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_175_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12688_ _03734_ _05950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_14427_ _00281_ net3 mod.u_cpu.rf_ram.memory\[474\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11639_ _05177_ _05234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_30_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08589__A1 _01496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_190_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12385__A2 _05726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_200_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14358_ _00212_ net3 mod.u_cpu.rf_ram.memory\[508\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_183_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10396__A1 _04389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_183_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13966__I _05801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_13309_ _06405_ _06406_ _06407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_144_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14289_ _00143_ net3 mod.u_cpu.rf_ram.memory\[543\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07651__I3 mod.u_cpu.rf_ram.memory\[299\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07964__I _01537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_237_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11196__I0 _04916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08436__S1 _02010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11486__I _03773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13885__A2 _06672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15546__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14420__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08850_ _02356_ mod.u_cpu.rf_ram.memory\[36\]\[1\] _03156_ _03157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_83_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07801_ _01701_ _02109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_131_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08761__A1 _03056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_257_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_242_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08781_ _02104_ _03068_ _03087_ _03088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_97_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_226_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_238_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11648__A1 _05239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07732_ _01444_ _02040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_66_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_226_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14570__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07316__A2 mod.u_cpu.rf_ram.memory\[484\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08513__A1 _01605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_211_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07663_ _01697_ mod.u_cpu.rf_ram.memory\[302\]\[0\] _01969_ _01970_ _01971_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_52_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_253_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10171__I1 _04111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_198_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09402_ _03637_ _03638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_198_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07594_ mod.u_cpu.rf_ram.memory\[352\]\[0\] mod.u_cpu.rf_ram.memory\[353\]\[0\] mod.u_cpu.rf_ram.memory\[354\]\[0\]
+ mod.u_cpu.rf_ram.memory\[355\]\[0\] _01841_ _01844_ _01902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_129_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_244_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09333_ _03578_ _03579_ _03580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__12073__A1 _05417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_205_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08744__B _01481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09264_ _03520_ _03521_ _03522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_138_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08215_ _02097_ _02523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_53_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09195_ mod.u_arbiter.i_wb_cpu_rdt\[23\] mod.u_arbiter.i_wb_cpu_dbus_dat\[20\] _03469_
+ _03470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_147_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_194_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15076__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08146_ _02453_ _02454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_146_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_193_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08077_ _01924_ _02385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_162_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_162_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_161_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13876__A2 _06837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_249_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_216_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14913__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14125__I0 _07041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_130_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08979_ mod.u_cpu.cpu.state.init_done _03284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_4825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_217_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11990_ _05464_ mod.u_cpu.rf_ram.memory\[559\]\[1\] _05475_ _05477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_4869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08504__A1 _02041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08355__I1 mod.u_cpu.rf_ram.memory\[489\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10941_ _04757_ _00487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_216_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_205_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_217_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13660_ _06671_ _06672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_44_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10872_ _04711_ _00464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_232_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__14053__A2 _06998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_12611_ _05891_ mod.u_cpu.rf_ram.memory\[153\]\[1\] _05897_ _05899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12064__A1 _05488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_243_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__12955__I _06131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_13591_ _06616_ _01278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_227_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__11111__I0 _04862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_231_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__13800__A2 _06772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_212_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15330_ _01106_ net3 mod.u_cpu.rf_ram.memory\[246\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_12542_ _05827_ mod.u_cpu.rf_ram.memory\[164\]\[0\] _05852_ _05853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__15419__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_185_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_212_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_185_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_196_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15261_ _00017_ net4 mod.u_arbiter.i_wb_cpu_rdt\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_40_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10475__I _04442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07491__A1 _01773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_200_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12473_ _05808_ _00968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_14212_ _03968_ _05120_ _07103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08115__S0 _02369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_200_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11424_ _05088_ _00639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_184_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15192_ _01045_ net3 mod.u_cpu.rf_ram.memory\[140\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_165_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09232__A2 _03493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15569__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14443__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14143_ _07060_ _01386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_126_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11355_ _05028_ mod.u_cpu.rf_ram.memory\[306\]\[0\] _05042_ _05043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_126_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07784__I _02091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10306_ _04163_ _04327_ _04328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08991__A1 _03260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14074_ _07016_ _01361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_125_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11286_ _04995_ _04996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_106_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11178__I0 _04916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13025_ _05535_ _06080_ _06187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_234_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10237_ _04276_ mod.u_cpu.rf_ram.memory\[483\]\[0\] _04278_ _04279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_79_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14593__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08743__A1 _02992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_239_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10168_ _03898_ _04230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_120_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14976_ _00830_ net3 mod.u_cpu.rf_ram.memory\[19\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10099_ _04179_ _00223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_82_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_208_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_212_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13927_ _06017_ _06903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_235_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11350__I0 _05028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_208_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_223_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13858_ _06435_ _06370_ _06436_ _06852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__14044__A2 _06989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_245_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12809_ mod.u_cpu.rf_ram.memory\[229\]\[1\] _06005_ _06027_ _06029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_16_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13789_ mod.u_arbiter.i_wb_cpu_rdt\[26\] _03449_ _03502_ _06790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07959__I _01614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_188_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15099__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_231_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15528_ _01299_ net3 mod.u_cpu.cpu.immdec.imm19_12_20\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08283__C _02080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07482__A1 _01740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15459_ _01233_ net3 mod.u_cpu.cpu.ctrl.o_ibus_adr\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_198_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_198_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08000_ _01716_ _02308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_15_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07609__I0 mod.u_cpu.rf_ram.memory\[312\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10369__A1 _04311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14936__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09951_ _01463_ _03722_ _04077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_131_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11169__I0 _04901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13858__A2 _06370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08902_ _02507_ _03208_ _03209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_103_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09882_ _03805_ _04003_ _04030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08734__A1 _02197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_253_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08833_ _01592_ _03130_ _03139_ _03140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__09782__I0 _03916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_100_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_170_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08764_ _02298_ _03070_ _03071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_73_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07715_ mod.u_cpu.rf_ram.memory\[269\]\[0\] _02023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__08458__C _02764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08695_ mod.u_cpu.rf_ram.memory\[197\]\[1\] _03002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_122_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14316__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07646_ _01918_ _01948_ _01953_ _01929_ _01954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_214_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_214_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12046__A1 _02226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13094__I0 _06230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07577_ _01874_ _01878_ _01883_ _01884_ _01885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_41_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_213_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09316_ _03563_ _03565_ _03566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13794__A1 _06726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09462__A2 _03687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14466__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_178_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07473__A1 _01779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09247_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[3\] _03507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_107_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_222_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_139_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_222_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09178_ _03460_ _00017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_147_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08129_ _02157_ _02436_ _02437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_108_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08812__I2 mod.u_cpu.rf_ram.memory\[14\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10080__I0 _04162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08973__A1 _03256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_257_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11140_ _04895_ _00548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_135_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__13849__A2 mod.u_arbiter.i_wb_cpu_rdt\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11071_ _04845_ _04848_ _04849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_5301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_1242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10907__I0 _04728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08725__A1 _02197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10022_ _04124_ _00201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_103_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_193_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11580__I0 _05194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_248_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14830_ _00684_ net3 mod.u_cpu.rf_ram.memory\[272\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_4633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3910 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_217_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3921 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_264_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3932 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08368__C _02109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_217_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3943 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14761_ _00615_ net3 mod.u_cpu.rf_ram.memory\[307\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11973_ _05465_ _00811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12285__A1 _05563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_217_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11332__I0 _05014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3954 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_16_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3965 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3976 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3987 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10924_ _04541_ _04746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_13712_ _06363_ _06712_ _06719_ _06135_ _06720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_72_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_264_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3998 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14692_ _00546_ net3 mod.u_cpu.rf_ram.memory\[341\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__15241__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07700__A2 _01996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14809__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12685__I _03944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13643_ _03390_ _06654_ _06137_ _06655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_10855_ _04640_ _04698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13085__I0 _06217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_260_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_198_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_72_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_201_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12588__A2 _05882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_13574_ mod.u_arbiter.i_wb_cpu_dbus_adr\[20\] mod.u_arbiter.i_wb_cpu_dbus_adr\[21\]
+ _06604_ _06607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_160_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10786_ _04238_ _04648_ _04652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09453__A2 _03679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__15391__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15313_ mod.u_scanchain_local.module_data_in\[69\] net4 net7 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_158_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12525_ _05164_ _04302_ _05842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_185_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_200_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14959__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12456_ mod.u_arbiter.i_wb_cpu_dbus_dat\[3\] _05793_ _05794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_15244_ _00019_ net4 mod.u_arbiter.i_wb_cpu_ack vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11399__I0 _05071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08831__C _02415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11407_ _05077_ _00633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_15175_ _01028_ net3 mod.u_cpu.rf_ram.memory\[147\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12126__S _05564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12387_ _05744_ _00946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_114_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14126_ _07049_ _01380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_11338_ _04795_ _05031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_181_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_141_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14057_ mod.u_arbiter.i_wb_cpu_rdt\[27\] _06998_ _07004_ mod.u_arbiter.i_wb_cpu_dbus_dat\[27\]
+ _07005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_11269_ _04982_ _04983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_122_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08716__A1 _01608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13008_ _06107_ mod.u_cpu.rf_ram.memory\[86\]\[0\] _06175_ _06176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_132_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_41_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08811__S1 _02386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14339__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14959_ _00813_ net3 mod.u_cpu.rf_ram.memory\[549\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_254_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07500_ mod.u_cpu.rf_ram.memory\[447\]\[0\] _01808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_223_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_208_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08480_ _02778_ _02779_ _02786_ _02007_ _02787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_90_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07431_ _01458_ _01739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__14489__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13076__I0 mod.u_cpu.rf_ram.memory\[105\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_223_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_211_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08327__S0 _02632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_250_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07362_ _01669_ _01670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__11626__I1 mod.u_cpu.rf_ram.memory\[262\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_189_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12823__I0 _06038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09101_ _03401_ _03402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_241_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_175_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07293_ _01536_ _01593_ _01600_ _01587_ _01601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_176_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09032_ _03334_ _03335_ _03336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_190_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_117_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11939__I _03780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15114__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09934_ _04054_ mod.u_cpu.rf_ram.memory\[528\]\[1\] _04063_ _04065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_89_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08707__A1 _02385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12503__A2 _03873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09755__I0 _03916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09865_ _04017_ _04018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_131_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_258_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_219_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10514__A1 _04168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11562__I0 _05178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09380__A1 _03616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08816_ mod.u_cpu.rf_ram.memory\[29\]\[1\] _03123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_133_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15264__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09796_ _03704_ _03938_ _03966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_85_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_227_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12267__A1 _05417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08747_ _02156_ mod.u_cpu.rf_ram.memory\[108\]\[1\] _03054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_2505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11314__I0 _05014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10117__I1 mod.u_cpu.rf_ram.memory\[500\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_260_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_199_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_183_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08678_ _02543_ _02981_ _02984_ _01632_ _02985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__10817__A2 _04669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13822__C _06753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_214_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_199_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07629_ _01643_ mod.u_cpu.rf_ram.memory\[308\]\[0\] _01936_ _01937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08916__C _02489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_242_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_199_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13067__I0 _06199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10640_ _04527_ _04389_ _04554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_146_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_194_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10571_ _04436_ _04507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_210_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_195_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12310_ _05691_ _00922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13519__A1 _06568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_195_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13290_ mod.u_arbiter.i_wb_cpu_rdt\[4\] mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat\[4\]
+ _06122_ _06388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_154_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12241_ _05604_ _05645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_182_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_206_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_218_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09319__I _03497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09994__I0 _04091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12172_ _05325_ _05576_ _05598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_123_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_107_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11123_ _04883_ mod.u_cpu.rf_ram.memory\[343\]\[0\] _04884_ _04885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_155_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15607__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11054_ _04827_ mod.u_cpu.rf_ram.memory\[353\]\[0\] _04835_ _04836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_89_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_190_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10005_ _03961_ _04087_ _04113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_249_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_5186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_77_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_114_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_265_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14813_ _00667_ net3 mod.u_cpu.rf_ram.memory\[281\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_4463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_114_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11305__I0 _05007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_149_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14631__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_236_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09123__A1 _03362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08557__S0 _01994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_14744_ _00598_ net3 mod.u_cpu.rf_ram.memory\[315\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_233_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11956_ _05450_ mod.u_cpu.rf_ram.memory\[218\]\[1\] _05453_ _05455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_189_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10907_ _04728_ mod.u_cpu.rf_ram.memory\[376\]\[0\] _04734_ _04735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_11887_ _05405_ _05406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_199_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_14675_ _00529_ net3 mod.u_cpu.rf_ram.memory\[350\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_60_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_232_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11608__I1 _05065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14781__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10838_ _04686_ _00455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_13626_ _06111_ _06112_ _06639_ _01290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_60_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_242_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13557_ _06597_ _01263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_10769_ _04496_ _04640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_201_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07532__S1 _01828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12508_ _05725_ _05831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_172_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13488_ _06537_ _06551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__15137__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14183__A1 _07026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15227_ _01080_ net3 mod.u_cpu.rf_ram.memory\[12\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_12_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12439_ _05778_ _00964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10663__I _04568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10044__I0 _04140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15158_ _01011_ net3 mod.u_cpu.rf_ram.memory\[155\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_99_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10744__A1 _04201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13974__I _06942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14109_ _07038_ _01374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_114_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15089_ _00943_ net3 mod.u_cpu.rf_ram.memory\[17\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_07980_ _02136_ _02287_ _02288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_99_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15287__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09737__I0 _03916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12497__A1 _05606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09362__A1 _03563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08289__B _02077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08796__S0 _02211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09650_ _03814_ _03851_ _03852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09362__B2 mod.u_arbiter.i_wb_cpu_dbus_adr\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08601_ _02323_ _02904_ _02907_ _01631_ _02908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__12249__A1 _05649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09581_ _03796_ _03797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_250_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_242_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_255_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08548__S0 _01802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08532_ _02059_ mod.u_cpu.rf_ram.memory\[300\]\[1\] _02839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_224_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13997__A1 mod.u_arbiter.i_wb_cpu_dbus_dat\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08463_ _01858_ _02769_ _02770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_169_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__13214__I _06320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13749__A1 _06335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07414_ _01633_ _01722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_211_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_196_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08394_ _02686_ _02690_ _02105_ _02700_ _02701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_51_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_148_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07345_ _01632_ _01639_ _01652_ _01618_ _01653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__07428__A1 _01446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_177_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07523__S1 _01830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_176_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07276_ _01528_ _01584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_178_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_164_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11669__I _05254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_164_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09015_ mod.u_cpu.cpu.state.o_cnt_r\[1\] _03320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_164_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__14504__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13921__A1 _06456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13921__B2 _06452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10735__A1 _04352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_215_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07600__A1 _01745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07882__I _02026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09917_ _04017_ _04054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_132_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_265_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14654__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10338__I1 mod.u_cpu.rf_ram.memory\[468\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_259_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09353__A1 _03415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10014__S _04119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_219_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09848_ _04006_ _00145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_74_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3003 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09803__S _03970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3014 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_247_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3025 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3036 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_218_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09779_ _03936_ mod.u_cpu.rf_ram.memory\[550\]\[1\] _03952_ _03954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_37_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3047 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_261_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3058 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_215_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11810_ _04808_ _03866_ _05352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_3069 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12790_ _06016_ _01077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_199_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09602__I _03757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_215_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_265_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_230_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11741_ _05249_ _05304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07667__A1 _01740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_2_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_199_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11463__A2 _04996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12660__A1 _05300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_230_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_199_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_214_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_202_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11672_ _05257_ _00718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_202_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14460_ _00314_ net3 mod.u_cpu.rf_ram.memory\[457\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08218__I _02084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_230_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07419__A1 _01705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10623_ _04537_ mod.u_cpu.rf_ram.memory\[423\]\[1\] _04540_ _04544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_13411_ _06502_ _01212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12963__I _06139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14391_ _00245_ net3 mod.u_cpu.rf_ram.memory\[492\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_161_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_224_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08711__S0 _01647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_183_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13342_ _06438_ _06390_ _06439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_167_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07514__S1 _01821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08092__A1 _02356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10554_ _04495_ _00362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_154_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10974__A1 _04227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14165__A1 _03670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13273_ _06322_ _06371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_170_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10485_ _04429_ _04450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_5_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09049__I _03352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15012_ _00866_ net3 mod.u_cpu.rf_ram.memory\[74\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12224_ _02330_ _05632_ _05633_ _00894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__13912__A1 _06471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10726__A1 _04611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09592__A1 _03374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12155_ _05586_ _00872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_9_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13727__C _06486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_257_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09719__I0 _03877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11106_ _04872_ _00537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_1_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12086_ _04973_ _05388_ _05540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07725__C _02007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10329__I1 mod.u_cpu.rf_ram.memory\[46\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_110_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11037_ _04824_ _00516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_49_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09895__A2 _04038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_224_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_237_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_218_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_206_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12988_ _06160_ _01131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_233_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_220_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08556__C _01812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14727_ _00581_ net3 mod.u_cpu.rf_ram.memory\[324\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_75_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11939_ _03780_ _05443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_206_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07122__A3 _01430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_177_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14658_ _00512_ net3 mod.u_cpu.rf_ram.memory\[358\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_177_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13609_ _03365_ _06625_ _06627_ _06628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_119_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_242_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_14589_ _00443_ net3 mod.u_cpu.rf_ram.memory\[393\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_159_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14527__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07130_ mod.u_cpu.rf_ram_if.rtrig0 _01439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__12954__A2 _06128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07830__A1 _02136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_145_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09958__I0 _04073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13903__A1 _03355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13918__B _06487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14677__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07963_ _02244_ mod.u_cpu.rf_ram.memory\[252\]\[0\] _02270_ _02271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_101_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_253_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_247_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07635__C _01768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08138__A2 _02419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09186__I1 mod.u_arbiter.i_wb_cpu_dbus_dat\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09702_ _03807_ _03892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_68_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07894_ _01779_ _02202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_114_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07207__I mod.u_cpu.raddr\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_261_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_229_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07897__A1 _02204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09633_ _03775_ _03838_ _03839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_56_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_216_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11952__I _03795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_243_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09564_ _03740_ mod.u_cpu.rf_ram.memory\[572\]\[0\] _03783_ _03784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_82_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08515_ _02759_ _02818_ _02821_ _02764_ _02822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_130_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_230_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_212_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09495_ _03374_ _03720_ _03721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_82_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15302__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_184_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_224_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08310__A2 mod.u_cpu.rf_ram.memory\[478\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08446_ _02730_ _02752_ _02753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_208_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_208_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_221_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_212_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13198__A2 _06304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08377_ _02656_ mod.u_cpu.rf_ram.memory\[428\]\[1\] _02684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__12245__I1 mod.u_cpu.rf_ram.memory\[196\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_183_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07877__I _01551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15452__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07328_ _01635_ _01636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_165_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08074__A1 _01483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_176_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07259_ _01495_ _01567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_30_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09949__I0 _04071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_180_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10270_ _04301_ _04302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_105_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_219_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11756__I0 _05304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10708__A1 _04168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08216__I3 mod.u_cpu.rf_ram.memory\[515\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09574__A1 _03758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08377__A2 mod.u_cpu.rf_ram.memory\[428\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_239_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_254_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08129__A2 _02436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09177__I1 mod.u_arbiter.i_wb_cpu_dbus_dat\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13960_ _03444_ _06917_ _06918_ _06931_ _06932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_47_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11133__A1 _04014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09877__A2 _04026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12911_ _06088_ mod.u_cpu.rf_ram.memory\[399\]\[0\] _06096_ _06097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_207_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12958__I _06134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_207_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13891_ _01426_ _06881_ _06800_ _01313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__12881__A1 _03968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11862__I _05387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_206_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_219_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15630_ _01401_ net3 mod.u_cpu.rf_ram.memory\[279\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12842_ _06038_ mod.u_cpu.rf_ram.memory\[123\]\[1\] _06049_ _06051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_185_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_226_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15561_ _01332_ net3 mod.u_arbiter.i_wb_cpu_dbus_dat\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07280__C _01587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12773_ _03734_ _06005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13830__B1 _06812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_215_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13830__C2 _06339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14512_ _00366_ net3 mod.u_cpu.rf_ram.memory\[431\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11724_ _05292_ _00735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_159_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_230_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15492_ _01263_ net3 mod.u_arbiter.i_wb_cpu_dbus_adr\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_203_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_120_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13189__A2 _06289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11655_ _05243_ mod.u_cpu.rf_ram.memory\[258\]\[0\] _05244_ _05245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_30_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14443_ _00297_ net3 mod.u_cpu.rf_ram.memory\[466\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_230_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10606_ _03733_ _04531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_11586_ _05198_ _00691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_200_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14374_ _00228_ net3 mod.u_cpu.rf_ram.memory\[500\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_10_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11995__I0 _05464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_183_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10798__I1 _04658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_183_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13325_ _06421_ _06422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_10537_ _04484_ _00356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_156_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10468_ _03991_ _04437_ _04438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_13256_ _06354_ mod.u_cpu.rf_ram.memory\[95\]\[1\] _06352_ _06355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_108_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_171_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11747__I0 _05304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08368__A2 mod.u_cpu.rf_ram.memory\[486\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12207_ _05621_ _00889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13361__A2 _06447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13187_ _06284_ _06294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_97_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10399_ mod.u_cpu.rf_ram.memory\[45\]\[1\] _04383_ _04390_ _04392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_151_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12138_ _05574_ _00867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_96_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_229_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09317__A1 _03415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12069_ _05521_ mod.u_cpu.rf_ram.memory\[63\]\[0\] _05528_ _05529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_226_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07879__A1 _02149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_253_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11675__A2 _05120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15325__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_38_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_225_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10722__I1 mod.u_cpu.rf_ram.memory\[406\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08540__A2 mod.u_cpu.rf_ram.memory\[292\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4090 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07194__I3 mod.u_cpu.rf_ram.memory\[451\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07974__S1 _02127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_53_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_241_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09242__I _03502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_212_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_206_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_206_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_209_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08300_ _02083_ _02598_ _02605_ _02606_ _02607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_178_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09280_ _03495_ _03535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_100_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15475__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08231_ _02120_ _02539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_159_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12309__S _05690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07697__I _01491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_147_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08056__A1 _02348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08162_ _02449_ _02452_ _02468_ _02469_ _02470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_140_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_158_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09253__B1 _03408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_140_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07113_ mod.u_cpu.cpu.branch_op _01422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_88_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_107_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08093_ _02352_ _02397_ _02400_ _02361_ _02401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_174_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_238_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_216_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_114_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_251_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10166__A2 _04227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08995_ _03280_ _03299_ _03300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11883__S _05402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09159__I1 mod.u_arbiter.i_wb_cpu_dbus_dat\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07946_ _02174_ _02248_ _02253_ _01766_ _02254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_87_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_205_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_214_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07877_ _01551_ _02185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_95_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_249_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09616_ _02513_ _03824_ _03825_ _00094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_141_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08196__C _02467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10298__I _03796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09547_ _03768_ _03749_ _03769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_231_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_212_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13603__S _06621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10477__I0 _04423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_212_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_196_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09478_ _01660_ _03703_ _03704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_70_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_211_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_200_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__14842__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08429_ _02534_ mod.u_cpu.rf_ram.memory\[404\]\[1\] _02735_ _02736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_138_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13415__I0 _06354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_184_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11123__S _04884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08047__A1 _02135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11440_ _05087_ mod.u_cpu.rf_ram.memory\[292\]\[1\] _05097_ _05099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_11_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09244__B1 _03497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09244__C2 mod.u_arbiter.i_wb_cpu_dbus_adr\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11371_ _05050_ mod.u_cpu.rf_ram.memory\[304\]\[1\] _05052_ _05054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_165_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08940__B _03246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13110_ _03960_ _06223_ _06242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_125_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10322_ _04338_ _00287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__14992__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14090_ _07026_ _07025_ _07027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_180_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13041_ _05606_ _06092_ _06197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13343__A2 _06418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10253_ _04289_ _00267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_140_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11354__A1 _04758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08231__I _02120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14222__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_182_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10184_ _04215_ mod.u_cpu.rf_ram.memory\[491\]\[1\] _04239_ _04241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07275__C _01582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15348__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10952__I1 mod.u_cpu.rf_ram.memory\[36\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08770__A2 _03069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14992_ _00846_ net3 mod.u_cpu.rf_ram.memory\[64\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12154__I0 _05575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_235_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12688__I _03734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13943_ _06912_ _06917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_93_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12854__A1 _06057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11901__I0 _05406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_207_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_262_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14372__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_235_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13874_ _06412_ _06834_ _06867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__15498__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_15613_ _01384_ net3 mod.u_cpu.rf_ram.memory\[115\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_74_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11409__A2 _05062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12825_ _03770_ _06030_ _06040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_76_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15544_ _01315_ net3 mod.u_cpu.rf_ram.memory\[112\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12756_ _05994_ _01065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_203_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08834__C _02380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10093__A1 _04044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11707_ _05265_ _05280_ _05281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_187_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15475_ _00005_ net3 mod.u_cpu.cpu.ctrl.pc_plus_4_cy_r vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12687_ _02370_ _05947_ _05949_ _01041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_129_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_204_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14426_ _00280_ net3 mod.u_cpu.rf_ram.memory\[474\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08038__A1 _02339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11638_ _05233_ _00708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08038__B2 _02345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07310__I _01551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08589__A2 mod.u_cpu.rf_ram.memory\[268\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14357_ _00211_ net3 mod.u_cpu.rf_ram.memory\[50\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_116_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_196_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11569_ _04066_ _05187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__11593__A1 _04930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10396__A2 _03896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_239_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13308_ _06374_ _06362_ _06406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_13_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_239_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14288_ _00142_ net3 mod.u_cpu.rf_ram.memory\[543\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_170_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10671__I _04574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13239_ _06343_ _01199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_171_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_258_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08141__I _02124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_151_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07800_ mod.u_cpu.rf_ram.memory\[168\]\[0\] mod.u_cpu.rf_ram.memory\[169\]\[0\] mod.u_cpu.rf_ram.memory\[170\]\[0\]
+ mod.u_cpu.rf_ram.memory\[171\]\[0\] _02106_ _02107_ _02108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_08780_ _01446_ _03077_ _03086_ _03087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_111_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13098__A1 _03950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14715__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07731_ _01485_ _02039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_266_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_226_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11648__A2 _03805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12845__A1 _01478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13893__I0 _06578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08297__B _02603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09710__A1 _03899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11208__S _04939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08513__A2 mod.u_cpu.rf_ram.memory\[348\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07662_ _01701_ _01970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_168_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10320__A2 _04336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09401_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[27\] mod.u_cpu.cpu.ctrl.o_ibus_adr\[26\] _03627_
+ _03637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__14865__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_179_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07593_ _01852_ _01892_ _01900_ _01677_ _01901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_213_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_213_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11007__I _04802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09332_ _03574_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[14\] _03560_ _03579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_80_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_240_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__12073__A2 _05388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_178_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_181_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09263_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[4\] mod.u_cpu.cpu.ctrl.o_ibus_adr\[3\] mod.u_cpu.cpu.ctrl.o_ibus_adr\[2\]
+ _03498_ _03521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_139_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_194_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_194_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08214_ _02039_ _02493_ _02521_ _02522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_09194_ _03451_ _03469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_222_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07220__I _01527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11959__I0 _05442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_193_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_147_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08145_ _01782_ _02453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_105_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_174_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08076_ mod.u_cpu.rf_ram.memory\[4\]\[0\] mod.u_cpu.rf_ram.memory\[5\]\[0\] mod.u_cpu.rf_ram.memory\[6\]\[0\]
+ mod.u_cpu.rf_ram.memory\[7\]\[0\] _02366_ _02383_ _02384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_162_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14245__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08051__I _01820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_102_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_248_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_88_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14395__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08978_ _01430_ mod.u_arbiter.i_wb_cpu_dbus_dat\[5\] mod.u_cpu.cpu.state.init_done
+ _03282_ _03283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_264_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07890__I _02197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_229_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15640__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_217_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07929_ mod.u_cpu.rf_ram.memory\[231\]\[0\] _02237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_112_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_217_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11118__S _04877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08504__A2 mod.u_cpu.rf_ram.memory\[324\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_244_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_217_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08060__S0 _02366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10940_ _04756_ mod.u_cpu.rf_ram.memory\[371\]\[1\] _04754_ _04757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_186_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10871_ _04695_ mod.u_cpu.rf_ram.memory\[382\]\[0\] _04710_ _04711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XPHY_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_12610_ _05898_ _01015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_71_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_197_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12064__A2 _05525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13261__A1 _06126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_13590_ mod.u_arbiter.i_wb_cpu_dbus_adr\[27\] mod.u_arbiter.i_wb_cpu_dbus_adr\[28\]
+ _06614_ _06616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_197_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08654__C _02141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12541_ _05367_ _05831_ _05852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_236_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_223_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_212_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_177_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15020__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08226__I _02216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15260_ _00016_ net4 mod.u_arbiter.i_wb_cpu_rdt\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12472_ _05807_ mod.u_cpu.rf_ram.memory\[419\]\[1\] _05804_ _05808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08115__S1 _02218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_14211_ _07102_ _01413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09768__A1 _03945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11423_ _05087_ mod.u_cpu.rf_ram.memory\[295\]\[1\] _05085_ _05088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_32_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15191_ _01044_ net3 mod.u_cpu.rf_ram.memory\[141\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_126_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_197_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11354_ _04758_ _05038_ _05042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_14142_ _07055_ mod.u_cpu.rf_ram.memory\[289\]\[1\] _07058_ _07060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_153_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08440__A1 _02143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_180_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15170__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10305_ _04302_ _04327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_153_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13316__A2 _06413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11285_ _04988_ _04995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_14073_ _06578_ mod.u_cpu.rf_ram.memory\[114\]\[0\] _07015_ _07016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_141_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14738__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12375__I0 _05731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11178__I1 mod.u_cpu.rf_ram.memory\[334\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10236_ _04277_ _04263_ _04278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_3_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_13024_ _06072_ _06186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_140_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11878__A2 _05398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09940__A1 _04044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08594__I2 mod.u_cpu.rf_ram.memory\[258\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09791__I1 mod.u_cpu.rf_ram.memory\[548\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10167_ _03896_ _04228_ _04229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_94_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_266_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14888__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14975_ _00829_ net3 mod.u_cpu.rf_ram.memory\[58\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10098_ _04178_ mod.u_cpu.rf_ram.memory\[503\]\[1\] _04174_ _04179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_130_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13926_ _02304_ _06901_ _06902_ _01327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_263_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13857_ _06487_ _06850_ _06851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_235_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_250_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_222_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12808_ _02234_ _06027_ _06028_ _01083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_90_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_204_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__13252__A1 _04984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_245_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_204_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13788_ mod.u_cpu.cpu.immdec.imm30_25\[1\] _06789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_204_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_231_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15527_ _01298_ net3 mod.u_cpu.cpu.immdec.imm19_12_20\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_206_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12739_ _02215_ _05982_ _05983_ _01059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_124_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_176_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15458_ _01232_ net3 mod.u_cpu.cpu.ctrl.o_ibus_adr\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__13004__A1 _01453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14268__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_191_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14409_ _00263_ net3 mod.u_cpu.rf_ram.memory\[483\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_102_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07609__I1 mod.u_cpu.rf_ram.memory\[313\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15513__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15389_ _01164_ net3 mod.u_cpu.rf_ram.memory\[103\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_117_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07975__I _02212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08431__A1 _02244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07865__S0 _02171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13307__A2 _06404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09950_ _04076_ _00177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08982__A2 mod.u_cpu.cpu.csr_d_sel vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_252_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11169__I1 mod.u_cpu.rf_ram.memory\[335\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08901_ mod.u_cpu.rf_ram.memory\[517\]\[1\] _03208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_106_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09881_ _04029_ _00155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_48_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08734__A2 _03040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09931__A1 _03873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08832_ _02150_ _03131_ _03138_ _02363_ _03139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_100_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_257_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08739__C _01695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08763_ mod.u_cpu.rf_ram.memory\[125\]\[1\] _03070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_111_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_211_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_211_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07714_ _01704_ _02022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_38_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08498__A1 _01875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08694_ _01560_ _03001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07215__I _01497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_253_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_226_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_199_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13618__I0 _06581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07645_ _01938_ mod.u_cpu.rf_ram.memory\[294\]\[0\] _01951_ _01952_ _01953_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_198_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_198_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15043__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12046__A2 _05512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07576_ _01630_ _01884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_41_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_241_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09315_ mod.u_arbiter.i_wb_cpu_dbus_adr\[13\] _03564_ _03565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_107_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13794__A2 _06407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14048__I _06963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_194_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09246_ _03493_ _03506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08670__A1 _02759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07473__A2 _01780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_182_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15193__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09177_ _03458_ mod.u_arbiter.i_wb_cpu_dbus_dat\[12\] _03459_ _03460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12791__I _05105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08128_ mod.u_cpu.rf_ram.memory\[45\]\[0\] _02436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_107_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_162_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08812__I3 mod.u_cpu.rf_ram.memory\[15\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08059_ _01524_ _02367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_162_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12357__I0 _05711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11070_ _04847_ _04848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_163_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_249_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_49_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10021_ _04115_ mod.u_cpu.rf_ram.memory\[514\]\[1\] _04122_ _04124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_118_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_49_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12232__S _05637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_88_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_102_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3900 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_3911 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_217_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13127__I _06252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3922 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_245_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14760_ _00614_ net3 mod.u_cpu.rf_ram.memory\[307\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3933 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11972_ _05464_ mod.u_cpu.rf_ram.memory\[217\]\[1\] _05462_ _05465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_3944 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12285__A2 _03859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3955 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07125__I mod.u_cpu.cpu.genblk3.csr.o_new_irq vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11332__I1 mod.u_cpu.rf_ram.memory\[310\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3966 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13711_ _06716_ _06718_ _06719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_186_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3977 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10923_ _04184_ _04713_ _04745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_72_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12966__I _01425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3988 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14691_ _00545_ net3 mod.u_cpu.rf_ram.memory\[342\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3999 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07161__A1 _01463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_232_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07161__B2 mod.u_cpu.cpu.immdec.imm24_20\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_189_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_204_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13642_ _03274_ _06653_ _06654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_16_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10854_ _04697_ _00460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_227_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10048__A1 _03752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__13785__A2 _06753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14410__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__15536__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_13573_ _06606_ _01270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_198_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10785_ _04651_ _00437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_185_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15312_ _00073_ net4 mod.u_scanchain_local.module_data_in\[69\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_12524_ _05841_ _00986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__10843__I0 _04682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_201_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08661__A1 _02450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_158_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_15243_ _00008_ net4 mod.timer_irq vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_157_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12455_ mod.u_arbiter.i_wb_cpu_dbus_dat\[2\] _03430_ mod.u_arbiter.i_wb_cpu_dbus_dat\[1\]
+ _05793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_184_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11399__I1 mod.u_cpu.rf_ram.memory\[2\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14560__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_184_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11406_ _05069_ mod.u_cpu.rf_ram.memory\[298\]\[1\] _05075_ _05077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_125_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_201_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15174_ _01027_ net3 mod.u_cpu.rf_ram.memory\[147\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08413__A1 _02539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12386_ _05731_ mod.u_cpu.rf_ram.memory\[177\]\[0\] _05743_ _05744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_125_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14125_ _07041_ mod.u_cpu.rf_ram.memory\[116\]\[1\] _07047_ _07049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_67_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11337_ _05030_ _00610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_141_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_141_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12348__I0 _05713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_193_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14056_ _06970_ _07004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09213__I0 mod.u_arbiter.i_wb_cpu_rdt\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_234_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11268_ _04194_ _04982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_140_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08716__A2 mod.u_cpu.rf_ram.memory\[228\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13238__S _06341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13007_ _03828_ _06080_ _06175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_140_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10219_ _04176_ _04266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_80_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07744__B _02051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11199_ _04918_ mod.u_cpu.rf_ram.memory\[330\]\[0\] _04934_ _04935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_239_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_228_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11720__A1 _05037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09515__I _03738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_208_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_208_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15066__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14958_ _00812_ net3 mod.u_cpu.rf_ram.memory\[549\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_82_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_235_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13909_ _06311_ _06861_ _06443_ _06647_ _06890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_63_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14889_ _00743_ net3 mod.u_cpu.rf_ram.memory\[23\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_251_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07430_ _01474_ _01738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_90_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_223_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__13076__I1 _05971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07361_ _01491_ _01669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08327__S1 _02633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_204_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13776__A2 _06714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_176_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09100_ _03385_ _03400_ _03401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_206_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14903__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08652__A1 _02136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07292_ _01505_ _01596_ _01599_ _01584_ _01600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_202_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_248_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09031_ _01435_ mod.u_cpu.cpu.decode.co_ebreak _01452_ _03335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_163_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08955__A2 _03259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11020__I _03949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12339__I0 _05711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09204__I0 mod.u_arbiter.i_wb_cpu_rdt\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09933_ _04064_ _00172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08530__S _02272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_217_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08707__A2 mod.u_cpu.rf_ram.memory\[236\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_219_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09864_ _03762_ _04017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15409__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08815_ mod.u_cpu.rf_ram.memory\[24\]\[1\] mod.u_cpu.rf_ram.memory\[25\]\[1\] mod.u_cpu.rf_ram.memory\[26\]\[1\]
+ mod.u_cpu.rf_ram.memory\[27\]\[1\] _02366_ _02367_ _03122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__08469__C _01887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09795_ _03965_ _00133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_227_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08746_ mod.u_cpu.rf_ram.memory\[109\]\[1\] _03053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_73_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14433__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08677_ _02462_ mod.u_cpu.rf_ram.memory\[214\]\[1\] _02983_ _02597_ _02984_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__15559__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07143__A1 _01431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_214_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07628_ _01934_ _01935_ _01936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10300__S _04323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08891__A1 _02479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_202_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11078__I0 _04843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13767__A2 _03391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07559_ _01503_ _01867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_224_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09435__A3 _03664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14583__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10825__I0 _04666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10570_ _04452_ _04506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_107_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08705__S _01807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08643__A1 _02116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09229_ _03410_ mod.u_scanchain_local.module_data_in\[38\] _03491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12227__S _05632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11131__S _04888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__12578__I0 _05869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12240_ _05644_ _00899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_182_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12171_ _05597_ _00877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_101_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_257_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11122_ _03879_ _04869_ _04884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_111_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_235_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11053_ _04285_ _04822_ _04835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_89_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15089__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08254__S0 _02560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_5143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10004_ _04112_ _00195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_5154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08379__C _02080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14812_ _00666_ net3 mod.u_cpu.rf_ram.memory\[281\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_4453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_264_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_218_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_217_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_123_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_205_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10269__A1 _04132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09123__A2 _03385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_233_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08557__S1 _02010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14743_ _00597_ net3 mod.u_cpu.rf_ram.memory\[316\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_123_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11955_ _05454_ _00804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_264_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07134__A1 mod.u_cpu.cpu.immdec.imm24_20\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_233_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_205_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10906_ _04732_ _04733_ _04734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_205_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08882__A1 _02457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_178_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14674_ _00528_ net3 mod.u_cpu.rf_ram.memory\[350\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_60_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14926__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11886_ _05404_ _05405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_162_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_260_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_220_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_220_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13625_ mod.u_cpu.cpu.genblk3.csr.timer_irq_r _06111_ _06639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_189_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10837_ _04682_ mod.u_cpu.rf_ram.memory\[387\]\[1\] _04684_ _04686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_164_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13556_ mod.u_arbiter.i_wb_cpu_dbus_adr\[12\] mod.u_arbiter.i_wb_cpu_dbus_adr\[13\]
+ _06594_ _06597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_186_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10768_ _04639_ _00432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_200_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12507_ _05830_ _00980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_146_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13487_ _06550_ _01240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_185_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10699_ _04593_ mod.u_cpu.rf_ram.memory\[410\]\[1\] _04591_ _04594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_172_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15226_ _01079_ net3 mod.u_cpu.rf_ram.memory\[12\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_218_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_195_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12438_ _05753_ mod.u_cpu.rf_ram.memory\[172\]\[0\] _05777_ _05778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_201_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11241__I0 _04952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15157_ _01010_ net3 mod.u_cpu.rf_ram.memory\[156\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_126_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12369_ _05732_ _04137_ _05733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_99_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14306__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10744__A2 _04623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11792__I1 _04954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14108_ _07028_ mod.u_cpu.rf_ram.memory\[117\]\[1\] _07036_ _07038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_99_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_15088_ _00942_ net3 mod.u_cpu.rf_ram.memory\[17\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_141_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11775__I _05106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14039_ _06990_ _06991_ _01351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_136_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input1_I io_in[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12741__I0 _05984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08796__S1 _02386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14456__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_256_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_228_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08600_ _02136_ mod.u_cpu.rf_ram.memory\[262\]\[1\] _02906_ _01504_ _02907_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_132_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_209_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_212_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09580_ _03795_ _03796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12600__S _05889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09181__S _03459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08548__S1 _01932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08531_ mod.u_cpu.rf_ram.memory\[301\]\[1\] _02838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_51_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08462_ mod.u_cpu.rf_ram.memory\[373\]\[1\] _02769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_51_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_247_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07676__A2 mod.u_cpu.rf_ram.memory\[276\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_211_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10680__A1 _04542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07413_ _01696_ _01699_ _01718_ _01720_ _01721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_250_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13749__A2 _03428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08393_ _02083_ _02691_ _02699_ _02606_ _02700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_149_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_259_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07344_ _01572_ _01642_ _01650_ _01651_ _01652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_177_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07275_ _01577_ mod.u_cpu.rf_ram.memory\[470\]\[0\] _01580_ _01582_ _01583_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__12047__S _05512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_164_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09014_ _03297_ _03298_ _03255_ _03318_ _03319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_191_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08324__I _02347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12185__A1 _05606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_191_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09976__I1 _03925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_191_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13921__A2 _06468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15231__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11932__A1 _03892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10735__A2 _04599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_254_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07600__A2 mod.u_cpu.rf_ram.memory\[358\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09916_ _04053_ _00166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_99_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08236__S0 _02507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13685__A1 _06694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_258_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_219_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_219_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09847_ _03999_ mod.u_cpu.rf_ram.memory\[542\]\[1\] _04004_ _04006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_86_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15381__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3004 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_246_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3015 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09778_ _03953_ _00128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3026 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14949__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3037 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3048 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11299__I0 _04978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3059 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08927__C _02505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_227_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08729_ _02632_ mod.u_cpu.rf_ram.memory\[246\]\[1\] _03035_ _01702_ _03036_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_2325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_215_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_265_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_215_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11999__A1 _02221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_199_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11740_ _05303_ _00740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_199_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10030__S _04129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08864__A1 _02456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_242_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_230_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07403__I _01710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_202_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11671_ _05243_ mod.u_cpu.rf_ram.memory\[250\]\[0\] _05256_ _05257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_144_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_230_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12799__I0 _06019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13410_ _06354_ mod.u_cpu.rf_ram.memory\[91\]\[1\] _06500_ _06502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_169_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10622_ _01760_ _04540_ _04543_ _00382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_14390_ _00244_ net3 mod.u_cpu.rf_ram.memory\[492\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_122_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_31_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_13341_ _06374_ _06438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08711__S1 _01732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_195_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10553_ _04486_ mod.u_cpu.rf_ram.memory\[433\]\[0\] _04494_ _04495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_6_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08092__A2 mod.u_cpu.rf_ram.memory\[30\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14329__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10974__A2 _04779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_183_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13272_ _06369_ _06370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08234__I _01688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10484_ _01803_ _04448_ _04449_ _00338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_15011_ _00865_ net3 mod.u_cpu.rf_ram.memory\[208\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12223_ _05581_ _05632_ _05633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_108_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13912__A2 _06823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_194_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12154_ _05575_ mod.u_cpu.rf_ram.memory\[206\]\[0\] _05585_ _05586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_29_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14479__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11105_ _04862_ mod.u_cpu.rf_ram.memory\[346\]\[1\] _04870_ _04872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_155_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10205__S _04256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12085_ _05520_ _05539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13676__A1 _06437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13676__B2 _06372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11036_ _04803_ mod.u_cpu.rf_ram.memory\[356\]\[0\] _04823_ _04824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_249_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_238_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_231_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_265_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13428__A1 _03371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_266_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_218_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10939__I _04719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12987_ _06158_ mod.u_cpu.cpu.genblk3.csr.mcause31 _06159_ _06160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_3571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13315__I _06412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14726_ _00580_ net3 mod.u_cpu.rf_ram.memory\[324\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11938_ _05412_ _05442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08855__A1 _03017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_261_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15104__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10662__A1 _03993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_232_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14657_ _00511_ net3 mod.u_cpu.rf_ram.memory\[35\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_221_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11869_ _05385_ mod.u_cpu.rf_ram.memory\[72\]\[0\] _05392_ _05393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_21_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13608_ _03381_ _06626_ _06627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_60_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_193_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08607__A1 _01481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13600__A1 _03713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14588_ _00442_ net3 mod.u_cpu.rf_ram.memory\[393\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_159_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_220_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_201_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_201_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13539_ _06587_ _01255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_199_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15254__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12167__A1 _05593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15209_ _01062_ net3 mod.u_cpu.rf_ram.memory\[219\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_160_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13903__A2 _06140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09032__A1 _03334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07983__I _01533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07962_ _02245_ _02269_ _02270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_102_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09701_ _03891_ _00113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_67_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07893_ _02198_ _02199_ _02200_ _02201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_67_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07346__A1 _01489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_228_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09632_ _03834_ _03837_ _03838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_216_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_255_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09563_ _03758_ _03782_ _03783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_83_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08514_ _02526_ _02819_ _02820_ _01501_ _02821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_252_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_212_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08846__A1 _02365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09494_ _01448_ _01454_ _03719_ _03720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_224_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_196_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08445_ mod.u_cpu.rf_ram.memory\[396\]\[1\] mod.u_cpu.rf_ram.memory\[397\]\[1\] mod.u_cpu.rf_ram.memory\[398\]\[1\]
+ mod.u_cpu.rf_ram.memory\[399\]\[1\] _02751_ _02748_ _02752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_251_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_260_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08376_ mod.u_cpu.rf_ram.memory\[429\]\[1\] _02683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_149_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14056__I _06970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07327_ _01634_ _01635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_104_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09271__A1 _03506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_178_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07258_ _01536_ _01555_ _01565_ _01552_ _01566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_87_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14621__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07189_ mod.u_cpu.raddr\[1\] _01497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09023__A1 _03306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_258_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10708__A2 _04599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11756__I1 mod.u_cpu.rf_ram.memory\[238\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09574__A2 _03791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10025__S _04126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13658__A1 _06667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14771__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_259_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_232_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12910_ _04913_ _04570_ _06096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_115_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_247_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13890_ _06704_ _06881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12881__A2 _06048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09613__I _03822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_261_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15127__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12841_ _06050_ _01094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_62_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07561__C _01631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_266_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14083__A1 _03865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13130__I0 mod.u_arbiter.i_wb_cpu_rdt\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15560_ _01331_ net3 mod.u_arbiter.i_wb_cpu_dbus_dat\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12772_ _06004_ _01071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08229__I _01747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09885__I0 _04018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_243_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14511_ _00365_ net3 mod.u_cpu.rf_ram.memory\[432\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_64_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11723_ _05287_ mod.u_cpu.rf_ram.memory\[243\]\[1\] _05290_ _05292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_214_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_203_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15491_ _01262_ net3 mod.u_arbiter.i_wb_cpu_dbus_adr\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15277__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14442_ _00296_ net3 mod.u_cpu.rf_ram.memory\[466\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_230_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11654_ _04831_ _05214_ _05244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_175_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_202_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12397__A1 _05581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08392__C _02196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10605_ _04530_ _00378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_155_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14373_ _00227_ net3 mod.u_cpu.rf_ram.memory\[501\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11585_ _05194_ mod.u_cpu.rf_ram.memory\[26\]\[1\] _05196_ _05198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_167_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_156_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13324_ _06064_ _06421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_128_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10536_ _04469_ mod.u_cpu.rf_ram.memory\[436\]\[0\] _04483_ _04484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12149__A1 _02181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13255_ _06236_ _06354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09014__A1 _03297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10467_ _04436_ _04437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_170_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12206_ _05609_ mod.u_cpu.rf_ram.memory\[200\]\[1\] _05619_ _05621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_123_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13186_ _06292_ _06293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_151_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08612__I1 mod.u_cpu.rf_ram.memory\[133\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10398_ _02436_ _04390_ _04391_ _00310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_124_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12137_ _05566_ mod.u_cpu.rf_ram.memory\[74\]\[1\] _05572_ _05574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_150_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09317__A2 mod.u_scanchain_local.module_data_in\[50\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12068_ _04294_ _04845_ _05528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_96_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11019_ _04811_ _00511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_38_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_237_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4080 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4091 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_234_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_127_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10635__A1 _04272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_221_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14709_ _00563_ net3 mod.u_cpu.rf_ram.memory\[333\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_233_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_205_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08230_ _02533_ mod.u_cpu.rf_ram.memory\[518\]\[0\] _02536_ _02537_ _02538_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_127_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_159_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14644__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08161_ _02143_ _02469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08056__A2 _02351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09253__A1 _03479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09253__B2 mod.u_arbiter.i_wb_cpu_dbus_adr\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07112_ mod.u_cpu.cpu.decode.opcode\[2\] _01421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08092_ _02356_ mod.u_cpu.rf_ram.memory\[30\]\[0\] _02399_ _02359_ _02400_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_119_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_162_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_256_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_161_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12325__S _05700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13888__B2 _06879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14794__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_255_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10410__I1 _04383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08994_ mod.u_cpu.cpu.bne_or_bge _03299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_130_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07945_ _02249_ mod.u_cpu.rf_ram.memory\[238\]\[0\] _02251_ _02252_ _02253_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_130_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07319__A1 _01577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12163__I1 _05468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_217_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07876_ _02174_ _02178_ _02183_ _02166_ _02184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_110_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09433__I mod.u_cpu.cpu.immdec.imm11_7\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_243_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09615_ _03775_ _03824_ _03825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_55_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09546_ _03701_ _03768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_71_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_225_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_221_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_93_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_197_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10477__I1 mod.u_cpu.rf_ram.memory\[446\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_262_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_212_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09477_ _01439_ _01494_ mod.u_cpu.raddr\[1\] _03703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_245_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_169_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08428_ _02526_ _02734_ _02735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_212_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12379__A1 _05293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__08047__A2 mod.u_cpu.rf_ram.memory\[68\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08359_ _01762_ _02666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09244__A1 _03496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11370_ _05053_ _00620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_166_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10321_ _04330_ mod.u_cpu.rf_ram.memory\[471\]\[1\] _04336_ _04338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_153_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13040_ _06196_ _01147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_180_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13343__A3 _06403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10252_ _04288_ mod.u_cpu.rf_ram.memory\[481\]\[1\] _04286_ _04289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_156_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_191_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07558__A1 _01864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10183_ _04240_ _00246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_79_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14991_ _00845_ net3 mod.u_cpu.rf_ram.memory\[63\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12303__A1 _05452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_232_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_208_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12154__I1 mod.u_cpu.rf_ram.memory\[206\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13942_ _06123_ _06906_ _06911_ _03431_ _06916_ _01329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_115_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14517__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_219_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_189_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_235_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13873_ _06739_ mod.u_arbiter.i_wb_cpu_rdt\[7\] _06865_ _06866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_47_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07291__C _01582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13103__I0 _06237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07730__A1 _01481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_235_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15612_ _01383_ net3 mod.u_cpu.rf_ram.memory\[115\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_90_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_216_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12824_ _06039_ _01088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_62_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_262_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_215_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__14667__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15543_ _01314_ net3 mod.u_cpu.rf_ram.memory\[112\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12755_ _05992_ mod.u_cpu.rf_ram.memory\[80\]\[0\] _05993_ _05994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_91_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_188_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07798__I _01672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_203_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11706_ _04994_ _05279_ _05280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10093__A2 _04174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15474_ _01248_ net3 mod.u_cpu.cpu.ctrl.o_ibus_adr\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_231_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_188_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12686_ _05948_ _05947_ _05949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_243_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_147_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_198_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11417__I0 _05069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14425_ _00279_ net3 mod.u_cpu.rf_ram.memory\[475\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11637_ _05222_ mod.u_cpu.rf_ram.memory\[260\]\[0\] _05232_ _05233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_128_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11042__A1 _04277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_196_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14356_ _00210_ net3 mod.u_cpu.rf_ram.memory\[50\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11568_ _05186_ _00685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_156_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_171_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11593__A2 _05191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13307_ _06368_ _06404_ _06405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_143_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10519_ _04251_ _03911_ _04473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_196_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14287_ _00141_ net3 mod.u_cpu.rf_ram.memory\[544\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11499_ _05114_ mod.u_cpu.rf_ram.memory\[283\]\[0\] _05140_ _05141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_196_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_196_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_226_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_13238_ _06276_ mod.u_cpu.rf_ram.memory\[94\]\[1\] _06341_ _06343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_108_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13590__I0 mod.u_arbiter.i_wb_cpu_dbus_adr\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_174_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13169_ _06277_ _01195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_111_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_211_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13098__A2 _06223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07730_ _01481_ _01817_ _02037_ _01469_ _02038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_66_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10156__I0 _04217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15442__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12845__A2 _06052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08297__C _02093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_225_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07661_ _01967_ _01968_ _01969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09710__A2 _03897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_168_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07721__A1 _02027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_214_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09400_ _03635_ _03632_ _03636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_241_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_207_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07592_ _01874_ _01896_ _01899_ _01884_ _01900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_81_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_207_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09331_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[16\] _03578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__15592__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09474__A1 _01418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09262_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[5\] _03520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_194_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_194_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_244_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08213_ _02506_ _02519_ _02520_ _02521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_21_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09193_ _03468_ _00025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_159_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12081__I0 _05521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08144_ mod.u_cpu.rf_ram.memory\[544\]\[0\] mod.u_cpu.rf_ram.memory\[545\]\[0\] mod.u_cpu.rf_ram.memory\[546\]\[0\]
+ mod.u_cpu.rf_ram.memory\[547\]\[0\] _02450_ _02451_ _02452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_88_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_174_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08760__C _02363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08075_ _01524_ _02383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_134_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12908__I0 _06086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_216_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_161_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11894__S _05409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12533__A1 _01775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_142_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_130_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_102_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08977_ mod.u_cpu.cpu.state.stage_two_req _03282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_4805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13089__A2 _06227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07928_ _02175_ mod.u_cpu.rf_ram.memory\[228\]\[0\] _02235_ _02236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_116_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_4849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_256_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07859_ _02155_ _02160_ _02165_ _02166_ _02167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__14038__A1 mod.u_arbiter.i_wb_cpu_rdt\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08060__S1 _02367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10870_ _04299_ _04709_ _04710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_147_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_244_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_232_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_231_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_188_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08935__C _02555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_213_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13797__B1 _06790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09529_ _03715_ _03753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_71_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__11134__S _04891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_262_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_197_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11272__A1 _04746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_12540_ _05851_ _00992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_213_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_213_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_185_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__07411__I _01550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_197_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_197_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_184_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12471_ _05806_ _05807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_229_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_14210_ mod.u_cpu.rf_ram.memory\[269\]\[1\] _06221_ _07100_ _07102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_11422_ _05031_ _05087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_184_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09768__A2 _03943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15190_ _01043_ net3 mod.u_cpu.rf_ram.memory\[141\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_177_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08670__C _01872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15315__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14141_ _07059_ _01385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_126_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11353_ _05041_ _00615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_125_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08291__I2 mod.u_cpu.rf_ram.memory\[450\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_4_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10304_ _04248_ _04326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08242__I _02156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14072_ _03858_ _07014_ _07015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11284_ _03769_ _04994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_180_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13023_ _06185_ _01141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12375__I1 mod.u_cpu.rf_ram.memory\[17\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14180__S _07083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10235_ _03968_ _04277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_133_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15465__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_266_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10166_ _04225_ _04227_ _04228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_126_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07951__A1 _02245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_266_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_254_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_248_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14974_ _00828_ net3 mod.u_cpu.rf_ram.memory\[58\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12827__A2 _06040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10097_ _04177_ _04178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_94_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_208_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_207_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_13925_ _06249_ _06901_ _06902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_78_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_208_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10012__I _03995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13856_ _06397_ _06292_ _06850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_130_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_228_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13751__C _06330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_204_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12807_ _05948_ _06027_ _06028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_188_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13787_ _06774_ _06787_ _06788_ _01302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_15_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10999_ _04797_ mod.u_cpu.rf_ram.memory\[362\]\[1\] _04793_ _04798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_43_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_206_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_241_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11263__A1 _04838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15526_ _01297_ net3 mod.u_cpu.cpu.immdec.imm19_12_20\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12738_ _05843_ _05982_ _05983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12460__B1 _05797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10310__I0 _04330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_176_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_203_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15457_ _01231_ net3 mod.u_cpu.cpu.ctrl.o_ibus_adr\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_175_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12669_ _05709_ _05937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11015__A1 _04808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14408_ _00262_ net3 mod.u_cpu.rf_ram.memory\[483\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_15_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_191_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15388_ _01163_ net3 mod.u_cpu.rf_ram.memory\[104\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_144_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14154__I _06063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14339_ _00193_ net3 mod.u_cpu.rf_ram.memory\[518\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_239_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07865__S1 _02172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12515__A1 _05759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08900_ mod.u_cpu.rf_ram.memory\[512\]\[1\] mod.u_cpu.rf_ram.memory\[513\]\[1\] mod.u_cpu.rf_ram.memory\[514\]\[1\]
+ mod.u_cpu.rf_ram.memory\[515\]\[1\] _02494_ _02495_ _03207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_258_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09880_ _04018_ mod.u_cpu.rf_ram.memory\[537\]\[1\] _04027_ _04029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12603__S _05893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08814__S0 _02391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10377__I0 _04363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08195__A1 _02461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08831_ _02405_ _03134_ _03137_ _02415_ _03138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_170_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14832__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_170_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08762_ mod.u_cpu.rf_ram.memory\[120\]\[1\] mod.u_cpu.rf_ram.memory\[121\]\[1\] mod.u_cpu.rf_ram.memory\[122\]\[1\]
+ mod.u_cpu.rf_ram.memory\[123\]\[1\] _02294_ _02295_ _03069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_111_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_226_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07713_ mod.u_cpu.rf_ram.memory\[264\]\[0\] mod.u_cpu.rf_ram.memory\[265\]\[0\] mod.u_cpu.rf_ram.memory\[266\]\[0\]
+ mod.u_cpu.rf_ram.memory\[267\]\[0\] _02020_ _01995_ _02021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_22_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_238_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08693_ mod.u_cpu.rf_ram.memory\[192\]\[1\] mod.u_cpu.rf_ram.memory\[193\]\[1\] mod.u_cpu.rf_ram.memory\[194\]\[1\]
+ mod.u_cpu.rf_ram.memory\[195\]\[1\] _01578_ _01714_ _03000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__08498__A2 mod.u_cpu.rf_ram.memory\[334\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_199_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07644_ _01782_ _01952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_54_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_214_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14982__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_213_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_207_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07575_ _01879_ mod.u_cpu.rf_ram.memory\[374\]\[0\] _01881_ _01882_ _01883_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_22_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_210_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09314_ _03486_ _03564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_210_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07231__I _01538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_194_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09245_ _03505_ _00042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__15338__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_181_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_210_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_194_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_193_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__12054__I0 _05518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_182_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09176_ _03451_ _03459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_194_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_257_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11688__I _05221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12754__A1 _03872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08127_ mod.u_cpu.rf_ram.memory\[40\]\[0\] mod.u_cpu.rf_ram.memory\[41\]\[0\] mod.u_cpu.rf_ram.memory\[42\]\[0\]
+ mod.u_cpu.rf_ram.memory\[43\]\[0\] _02151_ _02383_ _02435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__11801__I0 _05329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10604__I1 _04396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_162_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14362__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15488__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08058_ _02058_ _02366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_162_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12357__I1 mod.u_cpu.rf_ram.memory\[122\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_248_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07233__I0 mod.u_cpu.rf_ram.memory\[456\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10020_ _04123_ _00200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_5314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07834__C _02141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_264_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11129__S _04888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_236_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_102_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_217_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3901 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3912 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_263_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3923 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13852__B _06483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11971_ _05405_ _05464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3934 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09686__A1 _03878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08489__A2 _02788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_179_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3945 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3956 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13710_ _06694_ _06363_ _06717_ _06718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_3967 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10922_ _04744_ _00481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_260_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3978 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14690_ _00544_ net3 mod.u_cpu.rf_ram.memory\[342\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3989 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_229_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09621__I _03828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07161__A2 mod.u_cpu.cpu.immdec.imm19_12_20\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_229_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08665__C _01696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13641_ _03297_ mod.u_cpu.cpu.decode.opcode\[1\] _06652_ _06653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_72_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10853_ _04695_ mod.u_cpu.rf_ram.memory\[384\]\[0\] _04696_ _04697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_72_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__10048__A2 _04143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_198_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08237__I _02325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13572_ mod.u_arbiter.i_wb_cpu_dbus_adr\[19\] mod.u_arbiter.i_wb_cpu_dbus_adr\[20\]
+ _06604_ _06606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12293__I0 _05679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_201_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10784_ _04641_ mod.u_cpu.rf_ram.memory\[396\]\[1\] _04649_ _04651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08110__A1 _01592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__11799__S _05344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_15311_ _00072_ net4 mod.u_scanchain_local.module_data_in\[68\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_158_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12523_ _05837_ mod.u_cpu.rf_ram.memory\[166\]\[1\] _05839_ _05841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XPHY_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_200_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__14705__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15242_ _01095_ net3 mod.u_cpu.rf_ram.memory\[123\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_185_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12454_ _03281_ _05791_ _05792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_173_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12745__A1 _02199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11405_ _05076_ _00632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_166_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15173_ _01026_ net3 mod.u_cpu.rf_ram.memory\[148\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12385_ _05742_ _05726_ _05743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08413__A2 _02712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_193_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_236_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14124_ _07048_ _01379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_197_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11336_ _05028_ mod.u_cpu.rf_ram.memory\[30\]\[0\] _05029_ _05030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_153_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14855__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14055_ mod.u_arbiter.i_wb_cpu_dbus_dat\[28\] _07000_ _07003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_97_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11267_ _04981_ _00589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_141_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10359__I0 _04363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12423__S _05768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13006_ _06174_ _01135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_171_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10218_ _04265_ _00256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_67_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11198_ _04792_ _04926_ _04934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_121_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07924__A1 _01977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10149_ _01648_ _04213_ _04214_ _00238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_255_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_212_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13762__B _06421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14957_ _00811_ net3 mod.u_cpu.rf_ram.memory\[217\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_130_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_208_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_208_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08856__B _03162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13908_ _03681_ _06641_ _06887_ _06889_ _01322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_36_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08348__S _01709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14888_ _00742_ net3 mod.u_cpu.rf_ram.memory\[23\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_250_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__14235__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_0 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_223_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13839_ _06138_ _06834_ _06835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__09429__A1 _03417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13053__I _06204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08147__I _02454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07360_ _01662_ _01667_ _01668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_94_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08101__A1 _02316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15509_ _01280_ net3 mod.u_arbiter.i_wb_cpu_dbus_adr\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_149_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07291_ _01545_ mod.u_cpu.rf_ram.memory\[502\]\[0\] _01598_ _01582_ _01599_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__07986__I _01864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14385__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09179__S _03459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09030_ _03290_ _03334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_175_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15630__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_191_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_191_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_264_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13536__I0 mod.u_arbiter.i_wb_cpu_dbus_adr\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09932_ _04051_ mod.u_cpu.rf_ram.memory\[528\]\[0\] _04063_ _04064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_116_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_259_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09204__I1 mod.u_arbiter.i_wb_cpu_dbus_dat\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09706__I _03895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09863_ _04016_ _00150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07915__A1 _02066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_213_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08814_ _03117_ _03118_ _03119_ _03120_ _02391_ _01720_ _03121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_218_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15010__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09794_ _03964_ mod.u_cpu.rf_ram.memory\[548\]\[1\] _03962_ _03965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07226__I _01533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_245_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08745_ mod.u_cpu.rf_ram.memory\[110\]\[1\] mod.u_cpu.rf_ram.memory\[111\]\[1\] _01508_
+ _03052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_38_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11971__I _05405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_242_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_187_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08676_ _01705_ _02982_ _02983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_183_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10522__I0 _04467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08340__A1 _02559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07627_ mod.u_cpu.rf_ram.memory\[309\]\[0\] _01935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_1828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15160__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_241_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_198_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__14728__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08057__I _02347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07558_ _01864_ _01865_ _01866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_167_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07526__S0 _01832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12975__A1 _03389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_195_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09435__A4 _03665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_195_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10825__I1 mod.u_cpu.rf_ram.memory\[38\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07489_ _01779_ _01796_ _01797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07896__I _01993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12027__I0 _05501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09228_ _03485_ _03490_ _00039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_167_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_210_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_194_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14878__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_177_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09159_ mod.u_arbiter.i_wb_cpu_rdt\[9\] mod.u_arbiter.i_wb_cpu_dbus_dat\[6\] _03442_
+ _03448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_135_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12170_ mod.u_cpu.rf_ram.memory\[205\]\[1\] _05468_ _05595_ _05597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_68_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13527__I0 _06578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11121_ _04882_ _04883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_122_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_249_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11052_ _04834_ _00521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11002__I1 _04658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_95_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08254__S1 _02561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07906__A1 _02209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10003_ mod.u_cpu.rf_ram.memory\[517\]\[1\] _04111_ _04109_ _04112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_265_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_237_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_4410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10761__I0 _04622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07136__I _01444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14811_ _00665_ net3 mod.u_cpu.rf_ram.memory\[282\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__14258__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12977__I _03269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11881__I _05262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15503__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14742_ _00596_ net3 mod.u_cpu.rf_ram.memory\[316\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11954_ _05442_ mod.u_cpu.rf_ram.memory\[218\]\[0\] _05453_ _05454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_18_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_218_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_205_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_232_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10905_ _04708_ _04733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_14673_ _00527_ net3 mod.u_cpu.rf_ram.memory\[351\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11885_ _05105_ _05404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_233_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_13624_ _06638_ _01289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_242_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10836_ _04685_ _00454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_164_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_186_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13555_ _06596_ _01262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_199_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10767_ _04637_ mod.u_cpu.rf_ram.memory\[398\]\[0\] _04638_ _04639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09831__A1 _03754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12018__I0 _05470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12506_ _05822_ mod.u_cpu.rf_ram.memory\[16\]\[1\] _05828_ _05830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_157_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_13486_ _03610_ _06545_ _06546_ _03616_ _06550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_160_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10698_ _04578_ _04593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_139_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_199_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15225_ _01078_ net3 mod.u_cpu.rf_ram.memory\[130\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12437_ _05325_ _05767_ _05777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_138_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_201_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11121__I _04882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08398__A1 _02500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_201_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_172_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15156_ _01009_ net3 mod.u_cpu.rf_ram.memory\[156\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11241__I1 mod.u_cpu.rf_ram.memory\[324\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12368_ _03849_ _05732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_154_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14107_ _02326_ _07036_ _07037_ _01373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_126_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11319_ _05014_ mod.u_cpu.rf_ram.memory\[312\]\[1\] _05016_ _05018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_15087_ _00941_ net3 mod.u_cpu.rf_ram.memory\[499\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__15033__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_180_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12299_ _05684_ _00918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_113_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09347__B1 _03402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14038_ mod.u_arbiter.i_wb_cpu_rdt\[22\] _06987_ _06982_ mod.u_arbiter.i_wb_cpu_dbus_dat\[22\]
+ _06991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_234_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_228_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_228_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_132_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08570__A1 _01963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_227_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15183__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_209_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08530_ mod.u_cpu.rf_ram.memory\[302\]\[1\] mod.u_cpu.rf_ram.memory\[303\]\[1\] _02272_
+ _02837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_224_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11457__A1 _05110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08322__A1 _02609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07756__S0 _02022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_251_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08461_ mod.u_cpu.rf_ram.memory\[368\]\[1\] mod.u_cpu.rf_ram.memory\[369\]\[1\] mod.u_cpu.rf_ram.memory\[370\]\[1\]
+ mod.u_cpu.rf_ram.memory\[371\]\[1\] _01837_ _01838_ _02768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_224_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_223_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08873__A2 mod.u_cpu.rf_ram.memory\[556\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07412_ _01719_ _01720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__12257__I0 _05635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_196_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08392_ _02188_ _02695_ _02698_ _02196_ _02699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_177_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_177_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07343_ _01528_ _01651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07428__A3 _01735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12009__I0 _05484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_148_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07274_ _01581_ _01582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_176_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12709__A1 _05870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09013_ _01431_ _03305_ _03311_ _03317_ _03318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_192_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_191_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12185__A2 _05568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_258_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11932__A2 _05319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09915_ _04051_ mod.u_cpu.rf_ram.memory\[531\]\[0\] _04052_ _04053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09889__A1 _03945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14400__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08236__S1 _02543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13685__A2 _06398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15526__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_247_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09846_ _04005_ _00144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_63_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3005 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09777_ _03916_ mod.u_cpu.rf_ram.memory\[550\]\[0\] _03952_ _03953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_3016 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_234_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3027 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3038 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08728_ _02084_ _03034_ _03035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_3049 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14550__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_214_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07747__S0 _01893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11999__A2 _05481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08659_ mod.u_cpu.rf_ram.memory\[221\]\[1\] _02966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_27_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10120__A1 _03722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_261_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08864__A2 mod.u_cpu.rf_ram.memory\[548\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_199_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11670_ _04868_ _05255_ _05256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_199_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_230_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_224_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__12948__A1 _06122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10621_ _04542_ _04540_ _04543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_23_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13340_ _06436_ _06437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_139_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10552_ _04360_ _04487_ _04494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_128_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_259_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_211_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_13271_ _06367_ _06368_ _06369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_155_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10483_ _04439_ _04448_ _04449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__15056__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15010_ _00864_ net3 mod.u_cpu.rf_ram.memory\[208\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_136_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12222_ _05019_ _05631_ _05632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13373__A1 _06468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10187__A1 _04242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13912__A3 _06390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12153_ _05312_ _05568_ _05585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_64_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10982__I0 _04774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_190_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11104_ _04871_ _00536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09329__B1 _03555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12084_ _05538_ _00849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_2_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11035_ _04821_ _04822_ _04823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_77_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_209_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_264_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14201__B _06056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12487__I0 _05813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_206_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12986_ _06063_ _03335_ _03375_ _06159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_218_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_233_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14725_ _00579_ net3 mod.u_cpu.rf_ram.memory\[325\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_45_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11937_ _05441_ _00799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_205_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11116__I _04795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08855__A2 _03154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_260_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__12239__I0 mod.u_cpu.rf_ram.memory\[109\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2893 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11868_ _05343_ _05388_ _05392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_14656_ _00510_ net3 mod.u_cpu.rf_ram.memory\[35\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10662__A2 _04132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_159_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08853__C _02212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13607_ _03309_ _06625_ _06626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10819_ _04674_ _00448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_60_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11799_ _05342_ mod.u_cpu.rf_ram.memory\[232\]\[0\] _05344_ _05345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_207_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08607__A2 _02758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14587_ _00441_ net3 mod.u_cpu.rf_ram.memory\[394\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_158_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11611__A1 _04804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13538_ mod.u_arbiter.i_wb_cpu_dbus_adr\[4\] mod.u_arbiter.i_wb_cpu_dbus_adr\[5\]
+ _06584_ _06587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_173_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_158_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_174_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07291__A1 _01545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10891__S _04722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13469_ _06539_ _06540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_173_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12167__A2 _05594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15208_ _01061_ net3 mod.u_cpu.rf_ram.memory\[219\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_57_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09032__A2 _03335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14423__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15549__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15139_ _00992_ net3 mod.u_cpu.rf_ram.memory\[165\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_114_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07961_ mod.u_cpu.rf_ram.memory\[253\]\[0\] _02269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_99_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_229_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09700_ _03890_ mod.u_cpu.rf_ram.memory\[558\]\[1\] _03887_ _03891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_101_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_229_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_214_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07892_ _01517_ mod.u_cpu.rf_ram.memory\[218\]\[0\] _01714_ _02200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__14573__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12611__S _05897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13934__C _05800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_256_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08543__A1 _02216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09631_ _03836_ _03837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_68_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07932__C _02166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_216_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09562_ _03781_ _03782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_71_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07504__I _01787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08513_ _01605_ mod.u_cpu.rf_ram.memory\[348\]\[1\] _02820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_24_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09493_ _01448_ mod.u_cpu.cpu.immdec.imm11_7\[1\] _03719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08846__A2 _03152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_247_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_224_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_208_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08444_ _01919_ _02751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_168_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_225_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_211_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08375_ mod.u_cpu.rf_ram.memory\[430\]\[1\] mod.u_cpu.rf_ram.memory\[431\]\[1\] _02585_
+ _02682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_177_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__15079__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_220_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07326_ _01633_ _01634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_176_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07282__A1 _01486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07257_ _01505_ _01559_ _01564_ _01529_ _01565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_192_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_219_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07188_ _01495_ _01496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_145_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10169__A1 _04230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09023__A2 _03269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_191_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_173_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_254_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10964__I0 _04772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13107__A1 _02284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14916__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_160_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_266_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13658__A2 _06669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12705__I1 _05950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10716__I0 _04593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08534__A1 _02188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09829_ _03990_ _03991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_100_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12840_ _06035_ mod.u_cpu.rf_ram.memory\[123\]\[0\] _06049_ _06050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_2101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_262_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07414__I _01633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14083__A2 _07014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_104_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_265_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_215_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_161_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13860__B _06840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12771_ mod.u_cpu.rf_ram.memory\[133\]\[0\] _05971_ _06003_ _06004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_1411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_259_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_215_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_203_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_261_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_242_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11722_ _05291_ _00734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_14510_ _00364_ net3 mod.u_cpu.rf_ram.memory\[432\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_54_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15490_ _01261_ net3 mod.u_arbiter.i_wb_cpu_dbus_adr\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11653_ _05221_ _05243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14441_ _00295_ net3 mod.u_cpu.rf_ram.memory\[467\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_187_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_122_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10604_ mod.u_cpu.rf_ram.memory\[425\]\[0\] _04396_ _04529_ _04530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_211_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14372_ _00226_ net3 mod.u_cpu.rf_ram.memory\[501\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11584_ _05197_ _00690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_211_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14446__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_195_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13323_ mod.u_cpu.cpu.immdec.imm11_7\[1\] _06358_ _06420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_155_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10535_ _04189_ _04464_ _04483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_11_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_202_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13254_ _06353_ _01204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_109_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_129_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10466_ _04435_ _04436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09014__A2 _03298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13897__A2 _06881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12205_ _05620_ _00888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_124_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13185_ mod.u_arbiter.i_wb_cpu_rdt\[6\] mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat\[6\]
+ _06126_ _06292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_170_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14596__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10397_ _04230_ _04390_ _04391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_124_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09076__I _03377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_237_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08773__A1 _01682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12136_ _05573_ _00866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_111_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12067_ _05527_ _00843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13754__C _06065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_238_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08525__A1 _01874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11018_ _04797_ mod.u_cpu.rf_ram.memory\[35\]\[1\] _04809_ _04811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_133_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_265_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_238_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11380__I0 _05046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4070 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09025__B _03329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4081 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4092 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07324__I _01631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13770__B _03377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12969_ _03344_ _06144_ _06145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08384__S0 _02559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_261_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14708_ _00562_ net3 mod.u_cpu.rf_ram.memory\[333\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10635__A2 _04534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_244_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15221__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08583__C _02030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_178_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14639_ _00493_ net3 mod.u_cpu.rf_ram.memory\[368\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_221_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_220_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08160_ _02455_ _02460_ _02466_ _02467_ _02468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_193_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12632__I0 _05904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07111_ mod.u_cpu.cpu.decode.co_mem_word mod.u_cpu.cpu.bne_or_bge mod.u_cpu.cpu.csr_d_sel
+ _01420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_174_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15371__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08091_ _01823_ _02398_ _02399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_174_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14939__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09005__A2 _03309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11199__I0 _04918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13888__A2 _06640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_255_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08764__A1 _02298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09915__S _04052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08993_ _03253_ _03298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_87_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_173_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07944_ _01827_ _02252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_141_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13664__C _06134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09714__I _03766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09564__I0 _03740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08758__C _02359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_228_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07875_ _02179_ mod.u_cpu.rf_ram.memory\[206\]\[0\] _02182_ _02164_ _02183_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_21_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_217_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11371__I0 _05050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10323__A1 _04180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_229_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12140__I _05387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09614_ _03767_ _03823_ _03824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__14319__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_244_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__14065__A2 _06919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_209_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09545_ _03766_ _03767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_70_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_243_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13812__A2 _06772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_262_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_224_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_212_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_145_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09476_ _03701_ _03702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_52_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_184_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__09492__A2 _03717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_240_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14469__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08427_ mod.u_cpu.rf_ram.memory\[405\]\[1\] _02734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__10595__I _04522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_238_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08127__S0 _02151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12379__A2 _05726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08358_ _01991_ _02665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_196_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07255__A1 _01561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07309_ _01572_ _01611_ _01616_ _01584_ _01617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_221_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08289_ _02592_ _02595_ _02077_ _02596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_138_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10320_ _01579_ _04336_ _04337_ _00286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_109_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10251_ _04266_ _04288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_30_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12315__I _05694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10937__I0 _04753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14128__I0 _07043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08755__A1 _02532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10182_ _04217_ mod.u_cpu.rf_ram.memory\[491\]\[0\] _04239_ _04240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_120_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_266_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_14990_ _00844_ net3 mod.u_cpu.rf_ram.memory\[63\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_59_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_266_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08507__A1 _01540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13941_ _03431_ _06912_ _06915_ _06916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_120_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_247_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13872_ _03503_ mod.u_arbiter.i_wb_cpu_rdt\[23\] _06865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_75_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15244__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15611_ _01382_ net3 mod.u_cpu.rf_ram.memory\[118\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07730__A2 _01817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12823_ _06038_ mod.u_cpu.rf_ram.memory\[126\]\[1\] _06036_ _06039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_28_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14178__S _07083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_203_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_243_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15542_ _01313_ net3 mod.u_cpu.cpu.decode.op26 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12754_ _03872_ _05576_ _05993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_203_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11705_ _05262_ _05279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__15394__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12685_ _03944_ _05948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15473_ _01247_ net3 mod.u_cpu.cpu.ctrl.o_ibus_adr\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_230_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_203_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08118__S0 _02403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_203_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_202_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11636_ _04821_ _05214_ _05232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_14424_ _00278_ net3 mod.u_cpu.rf_ram.memory\[475\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_187_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_196_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07246__A1 _01489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11567_ _05178_ mod.u_cpu.rf_ram.memory\[272\]\[1\] _05184_ _05186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_200_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11042__A2 _04822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14355_ _00209_ net3 mod.u_cpu.rf_ram.memory\[510\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_155_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13306_ _06387_ _06404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_10518_ _04472_ _00349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_14286_ _00140_ net3 mod.u_cpu.rf_ram.memory\[544\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11498_ _05139_ _05125_ _05140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_109_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13237_ _06342_ _01198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_115_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_196_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10449_ _04423_ mod.u_cpu.rf_ram.memory\[450\]\[0\] _04424_ _04425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_152_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_156_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13168_ _06276_ mod.u_cpu.rf_ram.memory\[349\]\[1\] _06274_ _06277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__13590__I1 mod.u_arbiter.i_wb_cpu_dbus_adr\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12119_ _05550_ mod.u_cpu.rf_ram.memory\[210\]\[1\] _05560_ _05562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_135_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12161__S _05590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13099_ _06230_ mod.u_cpu.rf_ram.memory\[102\]\[0\] _06234_ _06235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_85_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_250_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09534__I _03757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_242_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10156__I1 mod.u_cpu.rf_ram.memory\[494\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07660_ mod.u_cpu.rf_ram.memory\[303\]\[0\] _01968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_168_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_226_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14047__A2 _06989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_226_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_207_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12058__A1 _05428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07591_ _01879_ mod.u_cpu.rf_ram.memory\[366\]\[0\] _01898_ _01867_ _01899_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_129_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12895__I _06018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11105__I0 _04862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14611__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_225_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_248_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_206_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07989__I _02091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09330_ _03546_ _03576_ _03577_ _00056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__11805__A1 _05348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_222_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09474__A2 _01645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_179_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_205_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09261_ _03506_ _03515_ _03519_ _00044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_60_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08212_ _01489_ _02520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_221_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14761__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_178_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09192_ mod.u_arbiter.i_wb_cpu_rdt\[22\] mod.u_arbiter.i_wb_cpu_dbus_dat\[19\] _03464_
+ _03468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_159_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_222_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08143_ _02152_ _02451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_119_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12230__A1 _05322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12081__I1 mod.u_cpu.rf_ram.memory\[212\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08985__A1 mod.u_cpu.cpu.state.o_cnt_r\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09709__I _03898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_174_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08074_ _01483_ _02336_ _02381_ _02382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_179_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15117__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_175_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10919__I0 _04728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08737__A1 _02084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07229__I _01515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13730__A1 _06456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12533__A2 _05846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12071__S _05528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15267__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08976_ _03251_ _03280_ _03281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_4806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_130_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08488__C _02096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_229_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07927_ _02157_ _02234_ _02235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_60_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12297__A1 _05139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07858_ _01765_ _02166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__14038__A2 _06987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14291__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07789_ _02096_ _02097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07899__I _01787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_225_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13797__B2 _06395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09528_ _03751_ _03752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XPHY_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_101_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_213_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_213_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09459_ _03395_ _03686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07476__A1 _01689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_212_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_197_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_212_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_200_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12470_ _05709_ _05806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_138_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11421_ _01950_ _05085_ _05086_ _00638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_177_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_193_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14140_ _07057_ mod.u_cpu.rf_ram.memory\[289\]\[0\] _07058_ _07059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08976__A1 _03251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11352_ _05032_ mod.u_cpu.rf_ram.memory\[307\]\[1\] _05039_ _05041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_165_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_137_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_193_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_153_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10303_ _04325_ _00281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08291__I3 mod.u_cpu.rf_ram.memory\[451\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_180_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14071_ _05630_ _07014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_11283_ _04993_ _00593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_180_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07139__I _01439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_193_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13022_ _06184_ mod.u_cpu.rf_ram.memory\[10\]\[1\] _06182_ _06185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08728__A1 _02084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_180_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10234_ _04248_ _04276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_105_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10535__A1 _04189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11583__I0 _05180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07400__A1 _01705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10165_ _04226_ _04227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_48_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14973_ _00827_ net3 mod.u_cpu.rf_ram.memory\[214\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10096_ _04176_ _04177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_208_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14634__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13924_ _04067_ _06030_ _06901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_208_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_63_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13855_ mod.u_arbiter.i_wb_cpu_rdt\[22\] mod.u_arbiter.i_wb_cpu_rdt\[6\] _06335_
+ _06849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_35_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_223_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_207_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_262_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_216_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12806_ _05226_ _05320_ _06027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__14784__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_204_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13786_ mod.u_cpu.cpu.immdec.imm30_25\[0\] _06774_ _06788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10998_ _04796_ _04797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09700__I0 _03890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_245_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15525_ _01296_ net3 mod.u_cpu.cpu.csr_imm vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_128_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11263__A2 _04969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12737_ _03865_ _05552_ _05982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12460__A1 _05792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12460__B2 mod.u_arbiter.i_wb_cpu_dbus_dat\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_231_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_204_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13540__S _06584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_203_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15456_ _01230_ net3 mod.u_cpu.cpu.ctrl.o_ibus_adr\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_163_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_12668_ _05936_ _01035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__14201__A2 _06151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10963__I _04719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14407_ _00261_ net3 mod.u_cpu.rf_ram.memory\[484\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11619_ _05208_ mod.u_cpu.rf_ram.memory\[263\]\[1\] _05218_ _05220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_156_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11015__A2 _03969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15387_ _01162_ net3 mod.u_cpu.rf_ram.memory\[104\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_204_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11060__S _04839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12599_ _05873_ _05891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09529__I _03715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10074__I0 _04157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_190_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13960__A1 _03444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14338_ _00192_ net3 mod.u_cpu.rf_ram.memory\[518\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_171_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10774__A1 _03723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14269_ _00123_ net3 mod.u_cpu.rf_ram.memory\[553\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_98_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08719__A1 _02751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13712__A1 _06363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12515__A2 _05835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10377__I1 mod.u_cpu.rf_ram.memory\[462\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08814__S1 _01720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_252_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08195__A2 mod.u_cpu.rf_ram.memory\[574\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09392__A1 _03496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08830_ _02410_ mod.u_cpu.rf_ram.memory\[22\]\[1\] _03136_ _01830_ _03137_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_170_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_258_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08761_ _03056_ _03058_ _02149_ _03067_ _03068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_39_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__13476__B1 _06540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_226_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_211_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07712_ _01993_ _02020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_66_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10203__I _03932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08692_ _02348_ _02998_ _02377_ _02999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_26_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09695__A2 _03886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07643_ _01949_ _01950_ _01951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13079__I0 mod.u_cpu.rf_ram.memory\[105\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_254_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_226_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_214_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07574_ _01749_ _01882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_181_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09313_ _03413_ _03563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_146_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12451__A1 _03700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08750__S0 _02106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09244_ _03496_ mod.u_scanchain_local.module_data_in\[39\] _03497_ _03504_ _03408_
+ mod.u_arbiter.i_wb_cpu_dbus_adr\[2\] _03505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai222_1
XFILLER_179_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_210_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_194_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12203__A1 _05343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09175_ mod.u_arbiter.i_wb_cpu_rdt\[15\] _03458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_222_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_194_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12066__S _05525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09439__I _03331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14507__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08126_ _02365_ _02426_ _02433_ _02168_ _02434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__12754__A2 _05576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_162_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08057_ _02347_ _02365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_123_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_162_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13703__A1 _06371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09758__I0 _03936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11565__I0 _05180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14657__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_163_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_102_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07933__A2 _02233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_233_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11317__I0 _05007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_188_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08959_ _03254_ mod.u_cpu.cpu.decode.opcode\[1\] _03263_ _03264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_248_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3902 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08011__C _02306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10113__I _03842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3913 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_99_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3924 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11970_ _02203_ _05462_ _05463_ _00810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_3935 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09686__A2 _03879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3946 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09902__I _04043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_217_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3957 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10921_ _04739_ mod.u_cpu.rf_ram.memory\[374\]\[1\] _04742_ _04744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_17_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3968 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_205_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3979 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11145__S _04898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13424__I _06510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_244_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13640_ _03297_ _03681_ _06652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10852_ _04290_ _04687_ _04696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_32_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_220_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_260_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_241_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_72_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_201_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10783_ _04650_ _00436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_13571_ _06605_ _01269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_164_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_213_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_185_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_15310_ _00071_ net4 mod.u_scanchain_local.module_data_in\[67\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_201_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12522_ _05840_ _00985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_40_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_184_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_201_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14195__A1 _07076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15241_ _01094_ net3 mod.u_cpu.rf_ram.memory\[123\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__13242__I0 _06273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12453_ _03289_ _03667_ _05791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_184_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_200_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10056__I0 _04148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11404_ _05071_ mod.u_cpu.rf_ram.memory\[298\]\[0\] _05075_ _05076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12745__A2 _05986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15432__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13942__A1 _06123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08253__I _02107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15172_ _01025_ net3 mod.u_cpu.rf_ram.memory\[148\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12384_ _03864_ _05742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_125_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_197_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_181_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11335_ _04196_ _03752_ _05029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_158_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14123_ _07043_ mod.u_cpu.rf_ram.memory\[116\]\[0\] _07047_ _07048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_21_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11266_ _04976_ mod.u_cpu.rf_ram.memory\[320\]\[1\] _04979_ _04981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_14054_ _07001_ _07002_ _01355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_106_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11556__I0 _05178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08016__I3 mod.u_cpu.rf_ram.memory\[115\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15582__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09374__A1 _03496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10217_ _04249_ mod.u_cpu.rf_ram.memory\[486\]\[0\] _04264_ _04265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__13170__A2 _03412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13005_ _06173_ mod.u_cpu.cpu.genblk3.csr.mcause3_0\[3\] _06163_ _06174_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_11197_ _04933_ _00567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_45_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11181__A1 _04643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_95_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07924__A2 _02187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_234_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10148_ _04186_ _04213_ _04214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_254_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14956_ _00810_ net3 mod.u_cpu.rf_ram.memory\[217\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10079_ _04163_ _04164_ _04165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_78_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08856__C _01891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09921__I0 _04051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13907_ _06647_ _06661_ _06682_ _06861_ _06888_ _06889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_236_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14887_ _00741_ net3 mod.u_cpu.rf_ram.memory\[240\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__13334__I _06133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13838_ _03331_ _03404_ _01424_ _03334_ _06834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_165_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_1 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_51_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_211_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_206_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_188_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12433__A1 _05642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13769_ _03670_ _03396_ _06771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_149_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08101__A2 mod.u_cpu.rf_ram.memory\[20\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_176_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08732__S0 _03001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_189_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15508_ _01279_ net3 mod.u_arbiter.i_wb_cpu_dbus_adr\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_07290_ _01561_ _01597_ _01598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_31_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08591__C _02764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15439_ _01214_ net3 mod.u_cpu.rf_ram.memory\[139\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_129_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09259__I _03517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13933__A1 _06153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_191_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08163__I _01688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09195__S _03469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09931_ _03873_ _04062_ _04063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11547__I0 _05159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13697__B1 _06450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09862_ _04001_ mod.u_cpu.rf_ram.memory\[53\]\[0\] _04015_ _04016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_252_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07915__A2 mod.u_cpu.rf_ram.memory\[214\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_259_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08813_ mod.u_cpu.rf_ram.memory\[8\]\[1\] mod.u_cpu.rf_ram.memory\[9\]\[1\] mod.u_cpu.rf_ram.memory\[10\]\[1\]
+ mod.u_cpu.rf_ram.memory\[11\]\[1\] _02171_ _02267_ _03120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09793_ _03889_ _03964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_133_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14110__A1 _03823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08744_ _02933_ _02965_ _01481_ _03050_ _03051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_227_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_27_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07679__A1 _01938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08675_ mod.u_cpu.rf_ram.memory\[215\]\[1\] _02982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_96_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_260_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_227_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15305__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_214_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_226_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_165_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_199_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07626_ _01710_ _01934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_148_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_183_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_242_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07557_ mod.u_cpu.rf_ram.memory\[383\]\[0\] _01865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_201_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_263_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08723__S0 _01647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_195_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07526__S1 _01833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_179_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__15455__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07488_ mod.u_cpu.rf_ram.memory\[439\]\[0\] _01796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_179_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_210_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09227_ _03371_ _03489_ _03490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07851__A1 _02157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_182_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_194_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13924__A1 _04067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09158_ _03446_ _03435_ _03447_ _00010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_147_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_194_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08109_ _02150_ _02404_ _02416_ _02363_ _02417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_181_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07603__A1 _01891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10108__I _04043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09089_ mod.u_cpu.cpu.state.o_cnt_r\[1\] _03388_ _03389_ mod.u_cpu.cpu.state.o_cnt_r\[2\]
+ _03390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_163_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_218_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11120_ _04620_ _04882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_122_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11538__I0 _05162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11051_ _04825_ mod.u_cpu.rf_ram.memory\[354\]\[1\] _04832_ _04834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_118_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_192_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_5101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_231_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_104_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_88_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10002_ _03928_ _04111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_118_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_190_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_191_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_236_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_249_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10761__I1 mod.u_cpu.rf_ram.memory\[3\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14810_ _00664_ net3 mod.u_cpu.rf_ram.memory\[282\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_4433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_218_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14741_ _00595_ net3 mod.u_cpu.rf_ram.memory\[317\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_218_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11953_ _05452_ _05423_ _05453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07580__C _01887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13154__I _06252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_229_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10904_ _03803_ _04732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_45_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14672_ _00526_ net3 mod.u_cpu.rf_ram.memory\[351\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11884_ _05403_ _00784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_45_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13623_ _06581_ mod.u_cpu.rf_ram.memory\[309\]\[1\] _06636_ _06638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_60_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12415__A1 _05588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10835_ _04679_ mod.u_cpu.rf_ram.memory\[387\]\[0\] _04684_ _04685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_220_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08692__B _02377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13090__S _06227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_13554_ mod.u_arbiter.i_wb_cpu_dbus_adr\[11\] mod.u_arbiter.i_wb_cpu_dbus_adr\[12\]
+ _06594_ _06596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_186_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09292__B1 _03536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10766_ _04218_ _04623_ _04638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_186_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14168__A1 _05790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12505_ _05829_ _00979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__14822__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12018__I1 mod.u_cpu.rf_ram.memory\[214\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_185_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13485_ _06549_ _01239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_10697_ _04592_ _00408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_186_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13915__A1 _05790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15224_ _01077_ net3 mod.u_cpu.rf_ram.memory\[130\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__13915__B2 _06465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12436_ _05776_ _00963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_173_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11777__I0 _05329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08398__A2 mod.u_cpu.rf_ram.memory\[436\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15155_ _01008_ net3 mod.u_cpu.rf_ram.memory\[157\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12367_ _05695_ _05731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__13757__C _06365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09807__I _03974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14972__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14106_ _07026_ _07036_ _07037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_11318_ _05017_ _00604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_141_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_259_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15086_ _00940_ net3 mod.u_cpu.rf_ram.memory\[499\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12298_ _05679_ mod.u_cpu.rf_ram.memory\[187\]\[0\] _05683_ _05684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__11529__I0 _05159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09347__A1 _03436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11249_ _04905_ _04969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_14037_ mod.u_arbiter.i_wb_cpu_dbus_dat\[23\] _06989_ _06990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09347__B2 mod.u_arbiter.i_wb_cpu_dbus_adr\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09028__B _03251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07327__I _01634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10201__I0 _04245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_132_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15328__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_255_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08570__A2 _02876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_250_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_247_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_242_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11457__A2 _03782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14939_ _00793_ net3 mod.u_cpu.rf_ram.memory\[223\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07490__C _01763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11701__I0 _05268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_208_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08460_ _01956_ _02766_ _01788_ _02767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__14352__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07756__S1 _02063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15478__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07411_ _01550_ _01719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_224_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08391_ _02191_ mod.u_cpu.rf_ram.memory\[422\]\[1\] _02697_ _02323_ _02698_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_56_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12609__S _05897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14096__S _07030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11513__S _05150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07342_ _01643_ mod.u_cpu.rf_ram.memory\[494\]\[0\] _01649_ _01615_ _01650_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_204_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12957__A2 _06133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10968__A1 _04775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14159__A1 _06153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07273_ _01523_ _01581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_177_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09012_ _03312_ _03287_ _03314_ _03315_ _03316_ _03317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__12709__A2 _04668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13906__A1 _06065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09918__S _04052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_191_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_191_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10440__I0 _04410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09717__I _03904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_219_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_219_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09914_ _03851_ _04038_ _04052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_217_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12193__I0 _05605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09889__A2 _04034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08010__A1 _02303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09845_ _04001_ mod.u_cpu.rf_ram.memory\[542\]\[0\] _04004_ _04005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_112_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_218_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09776_ _03948_ _03951_ _03952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_3006 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3017 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3028 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3039 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_227_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08727_ mod.u_cpu.rf_ram.memory\[247\]\[1\] _03034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_2305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_261_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_215_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13842__B1 _06837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_187_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07747__S1 _02054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_187_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08658_ _02944_ _02964_ _01738_ _02965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_42_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_226_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_215_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_241_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_230_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_215_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07609_ mod.u_cpu.rf_ram.memory\[312\]\[0\] mod.u_cpu.rf_ram.memory\[313\]\[0\] mod.u_cpu.rf_ram.memory\[314\]\[0\]
+ mod.u_cpu.rf_ram.memory\[315\]\[0\] _01774_ _01916_ _01917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_183_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14845__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_187_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_202_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08589_ _01496_ mod.u_cpu.rf_ram.memory\[268\]\[1\] _02896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_144_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11423__S _05085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12948__A2 _06123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10620_ _04541_ _04542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_41_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09813__A2 _03966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_195_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10551_ _04493_ _00361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_168_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_183_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14995__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13270_ _06120_ _06368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_10482_ _04307_ _04447_ _04448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_202_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13373__A2 _06403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12221_ _05630_ _05631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_204_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_135_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13912__A4 _06660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11384__A1 _03892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_194_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12152_ _05584_ _00871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_191_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_155_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__14225__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07575__C _01882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11103_ _04864_ mod.u_cpu.rf_ram.memory\[346\]\[0\] _04870_ _04871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_162_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10982__I1 mod.u_cpu.rf_ram.memory\[364\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09329__A1 _03554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12083_ _05533_ mod.u_cpu.rf_ram.memory\[212\]\[1\] _05536_ _05538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_78_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11034_ _04703_ _04822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08001__A1 _02283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_265_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_237_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13085__S _06224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14375__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_253_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15620__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_224_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12636__A1 _05535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12985_ _06113_ _03370_ _06158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_4296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14724_ _00578_ net3 mod.u_cpu.rf_ram.memory\[325\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11936_ mod.u_cpu.rf_ram.memory\[169\]\[1\] _05230_ _05439_ _05441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_3584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_127_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_221_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_206_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_178_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14655_ _00509_ net3 mod.u_cpu.rf_ram.memory\[360\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12239__I1 _05617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11867_ _05391_ _00779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_162_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2894 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_220_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08068__A1 _02352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13606_ _01429_ _03307_ _03315_ _06625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__13061__A1 _02353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10818_ _04663_ mod.u_cpu.rf_ram.memory\[390\]\[0\] _04673_ _04674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_198_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14586_ _00440_ net3 mod.u_cpu.rf_ram.memory\[394\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11798_ _05343_ _05335_ _05344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_186_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07610__I _01750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07815__A1 _01670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13537_ _06586_ _01254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_203_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_146_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10749_ _04627_ _00425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_174_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15000__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_174_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_199_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07291__A2 mod.u_cpu.rf_ram.memory\[502\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13468_ _06512_ _06539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_174_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_199_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_15207_ _01060_ net3 mod.u_cpu.rf_ram.memory\[209\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_126_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12419_ mod.u_cpu.rf_ram.memory\[489\]\[1\] _05765_ _05763_ _05766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_173_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13399_ _06310_ _06493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_99_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08441__I _01762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15138_ _00991_ net3 mod.u_cpu.rf_ram.memory\[165\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_142_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08240__A1 _02509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15150__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_141_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07960_ mod.u_cpu.rf_ram.memory\[248\]\[0\] mod.u_cpu.rf_ram.memory\[249\]\[0\] mod.u_cpu.rf_ram.memory\[250\]\[0\]
+ mod.u_cpu.rf_ram.memory\[251\]\[0\] _02266_ _02267_ _02268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_15069_ _00923_ net3 mod.u_cpu.rf_ram.memory\[185\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_114_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12175__I0 _05583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14718__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12898__I _06072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07891_ mod.u_cpu.rf_ram.memory\[219\]\[0\] _02199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__11922__I0 _05426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08543__A2 mod.u_cpu.rf_ram.memory\[294\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09630_ _03835_ _03836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_68_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09272__I _03488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_209_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09561_ _03780_ _03781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_23_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_243_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__14868__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08512_ mod.u_cpu.rf_ram.memory\[349\]\[1\] _02819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09492_ _03716_ _03717_ _03718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_64_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_223_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_212_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08443_ _01680_ _02749_ _02750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_169_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_212_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08374_ _02148_ _02680_ _02681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_23_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_225_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07520__I _01827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07325_ _01494_ _01633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07806__A1 _02111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07256_ _01545_ mod.u_cpu.rf_ram.memory\[478\]\[0\] _01563_ _01525_ _01564_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_192_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14248__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11977__I _05229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_178_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07187_ _01494_ _01495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_180_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10169__A2 _04229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08082__I1 mod.u_cpu.rf_ram.memory\[9\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_191_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13107__A2 _06239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_191_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14398__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12802__S _06024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_232_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_235_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15643__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_247_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_219_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11913__I0 _05413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08534__A2 _02837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09828_ _03749_ _03818_ _03990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_86_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_235_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_207_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_206_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09759_ _03937_ _00125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_64_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13633__S _03503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10121__I _04194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08298__A1 _02487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12770_ _04955_ _05952_ _06003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_64_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11721_ _05289_ mod.u_cpu.rf_ram.memory\[243\]\[0\] _05290_ _05291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_199_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13418__I0 _06351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_202_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_203_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11153__S _04902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15023__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14440_ _00294_ net3 mod.u_cpu.rf_ram.memory\[467\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11652_ _05242_ _00713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_187_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07430__I _01474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10603_ _04527_ _04528_ _04529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_128_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14371_ _00225_ net3 mod.u_cpu.rf_ram.memory\[502\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11583_ _05180_ mod.u_cpu.rf_ram.memory\[26\]\[0\] _05196_ _05197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_122_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13322_ _03664_ _06416_ _06339_ _06418_ _06419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_10_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10534_ _04482_ _00355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11887__I _05405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_196_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15173__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13253_ _06351_ mod.u_cpu.rf_ram.memory\[95\]\[0\] _06352_ _06353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_10465_ _03755_ _04132_ _04435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_170_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12204_ _05605_ mod.u_cpu.rf_ram.memory\[200\]\[0\] _05619_ _05620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_136_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10404__I0 _04387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08222__A1 _02528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13184_ _05783_ mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat\[5\] _06290_ _06291_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_151_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10396_ _04389_ _03896_ _04390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_151_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12135_ _05559_ mod.u_cpu.rf_ram.memory\[74\]\[0\] _05572_ _05573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_123_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12066_ _05518_ mod.u_cpu.rf_ram.memory\[29\]\[1\] _05525_ _05527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12857__A1 _01464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08525__A2 _02828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11017_ _04810_ _00510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08081__S0 _02266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07584__I0 mod.u_cpu.rf_ram.memory\[360\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11380__I1 mod.u_cpu.rf_ram.memory\[302\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4060 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_225_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4071 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4082 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11127__I _04847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4093 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_252_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08289__A1 _02592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_206_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13282__A1 _06328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_12968_ _06142_ _06143_ _06144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_248_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_206_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_205_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14707_ _00561_ net3 mod.u_cpu.rf_ram.memory\[334\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_73_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_221_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11919_ _05428_ _05423_ _05429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08384__S1 _02155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11063__S _04839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12899_ _03985_ _06048_ _06089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_178_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14638_ _00492_ net3 mod.u_cpu.rf_ram.memory\[368\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_21_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1990 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_147_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15516__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14569_ _00423_ net3 mod.u_cpu.rf_ram.memory\[403\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08836__I0 mod.u_cpu.rf_ram.memory\[48\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12632__I1 mod.u_cpu.rf_ram.memory\[14\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07110_ _01418_ mod.u_cpu.cpu.csr_imm _01419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_53_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08090_ mod.u_cpu.rf_ram.memory\[31\]\[0\] _02398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_158_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11797__I _03931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_174_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14540__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08171__I _01925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_251_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08992_ _03251_ _03297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_173_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_229_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07943_ _02180_ _02250_ _02251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_214_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12848__A1 _06052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14690__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_256_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09564__I1 mod.u_cpu.rf_ram.memory\[572\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_60_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12421__I _05725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_229_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_205_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07874_ _02180_ _02181_ _02182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_151_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_229_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_214_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09613_ _03822_ _03823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_3_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_249_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__15046__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09544_ _03756_ _03766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_37_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12320__I0 _05692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_212_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12069__S _05528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09475_ _01500_ _03700_ _03701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_224_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_197_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08426_ mod.u_cpu.rf_ram.memory\[400\]\[1\] mod.u_cpu.rf_ram.memory\[401\]\[1\] mod.u_cpu.rf_ram.memory\[402\]\[1\]
+ mod.u_cpu.rf_ram.memory\[403\]\[1\] _02688_ _02475_ _02733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_52_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10882__I0 _04695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13025__A1 _05535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_211_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__14073__I0 _06578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_200_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15196__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08127__S1 _02383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08357_ _01890_ _02664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_260_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07308_ _01577_ mod.u_cpu.rf_ram.memory\[510\]\[0\] _01613_ _01615_ _01616_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_165_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08288_ mod.u_cpu.rf_ram.memory\[456\]\[1\] mod.u_cpu.rf_ram.memory\[457\]\[1\] mod.u_cpu.rf_ram.memory\[458\]\[1\]
+ mod.u_cpu.rf_ram.memory\[459\]\[1\] _02593_ _02594_ _02595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_192_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_192_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13328__A2 _06304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07239_ _01520_ _01546_ _01547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_180_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10250_ _04287_ _00266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_180_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_145_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09952__A1 _03896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08014__C _02321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10181_ _04238_ _04234_ _04239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_160_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_266_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_160_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__12839__A1 _05888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13427__I _06513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08507__A2 mod.u_cpu.rf_ram.memory\[326\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09704__A1 _03702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13940_ _03434_ _06912_ _06914_ _06915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_87_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_235_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13871_ _06840_ _06859_ _06860_ _06863_ _06864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_207_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_262_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15610_ _01381_ net3 mod.u_cpu.rf_ram.memory\[118\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_75_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12822_ _06018_ _06038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_234_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_216_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_215_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_231_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_15541_ _01312_ net3 mod.u_cpu.cpu.immdec.imm24_20\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_128_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14413__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15539__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12753_ _05962_ _05992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_203_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11704_ _05278_ _00729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10873__I0 _04698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_188_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15472_ _01246_ net3 mod.u_cpu.cpu.ctrl.o_ibus_adr\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12684_ _03895_ _05589_ _05947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_70_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07160__I _01468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08118__S1 _02383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14423_ _00277_ net3 mod.u_cpu.rf_ram.memory\[476\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_175_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11635_ _05231_ _00707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_204_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14563__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14354_ _00208_ net3 mod.u_cpu.rf_ram.memory\[510\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08443__A1 _01680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11566_ _05185_ _00684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_129_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_171_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13305_ _06402_ _06403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_196_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10517_ _04467_ mod.u_cpu.rf_ram.memory\[440\]\[1\] _04470_ _04472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_14285_ _00139_ net3 mod.u_cpu.rf_ram.memory\[545\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_7_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11497_ _03789_ _05139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_100_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_171_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13236_ _06273_ mod.u_cpu.rf_ram.memory\[94\]\[0\] _06341_ _06342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_10448_ _04281_ _04407_ _04424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_124_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13538__S _06584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_237_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09794__I1 mod.u_cpu.rf_ram.memory\[548\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13167_ _06236_ _06276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_174_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10379_ _03894_ _04377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_124_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_258_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12118_ _05561_ _00860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_215_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13098_ _03950_ _06223_ _06234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_111_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13337__I _06125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_238_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12241__I _05604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__15069__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12049_ _03770_ _05515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_266_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_266_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_226_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07335__I _01604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_265_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07590_ _01663_ _01897_ _01898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_253_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12058__A2 _03878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_207_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_222_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_209_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_244_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_222_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09260_ _03516_ mod.u_scanchain_local.module_data_in\[41\] _03518_ mod.u_arbiter.i_wb_cpu_dbus_adr\[4\]
+ _03519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__13007__A1 _03828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14906__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08682__A1 _02477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_179_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08211_ _02471_ _02508_ _02517_ _02518_ _02519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_09191_ _03467_ _00024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_159_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12617__S _05901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_140_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08142_ _02209_ _02450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_147_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12230__A2 _05637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08073_ _02337_ _02346_ _02379_ _02380_ _02381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_175_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_255_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10919__I1 mod.u_cpu.rf_ram.memory\[374\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08737__A2 _03043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13730__A2 _06725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09725__I _03910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08769__C _02308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_102_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08975_ mod.u_cpu.cpu.decode.co_mem_word _03280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_9_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_257_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07926_ mod.u_cpu.rf_ram.memory\[229\]\[0\] _02234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_4829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_130_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_60_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12297__A2 _05668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09661__S _03860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13494__B2 _03635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14436__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07857_ _02161_ mod.u_cpu.rf_ram.memory\[198\]\[0\] _02163_ _02164_ _02165_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__07173__A1 _01478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_244_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08785__B _01720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_216_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__13246__A1 _03781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07788_ _01686_ _02096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_147_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_213_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_262_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09527_ _03750_ _03751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_240_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__14586__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08673__A1 _02202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09458_ mod.u_cpu.cpu.bufreg.c_r _03684_ _03685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_52_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07476__A2 mod.u_cpu.rf_ram.memory\[430\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_227_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08409_ mod.u_cpu.rf_ram.memory\[447\]\[1\] _02716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09389_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[25\] _03626_ _03627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_196_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_200_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11420_ _05022_ _05085_ _05086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_123_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_137_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08815__I3 mod.u_cpu.rf_ram.memory\[27\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11280__I0 _04978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11351_ _05040_ _00614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_138_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_197_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08025__B _02332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10302_ _04313_ mod.u_cpu.rf_ram.memory\[474\]\[1\] _04323_ _04325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_14070_ _03483_ _06911_ _06919_ _07012_ _07013_ _01360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_3_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11282_ _04976_ mod.u_cpu.rf_ram.memory\[318\]\[1\] _04991_ _04993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09925__A1 _04013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13021_ _06104_ _06184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_10233_ _04275_ _00261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_69_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_234_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15211__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10164_ _03992_ _04134_ _04226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_79_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14972_ _00826_ net3 mod.u_cpu.rf_ram.memory\[214\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10095_ _03761_ _04176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08036__S0 _01636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_266_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_247_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07155__I _01463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10299__A1 _04322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13923_ _06641_ _06899_ _06900_ _01326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_130_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07164__A1 _01462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15361__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_263_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11606__S _05211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13854_ _06847_ _06848_ _01309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_34_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_235_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14929__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_235_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12805_ _06026_ _01082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_90_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13785_ mod.u_cpu.cpu.immdec.imm30_25\[1\] _06753_ _06786_ _06787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_50_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10997_ _04795_ _04796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_245_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15524_ _01295_ net3 mod.u_cpu.cpu.immdec.imm19_12_20\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_16_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09700__I1 mod.u_cpu.rf_ram.memory\[558\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12736_ _05981_ _01058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08664__A1 _02566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_230_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10471__A1 _01808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15455_ _01229_ net3 mod.u_cpu.cpu.ctrl.o_ibus_adr\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12667_ _05934_ mod.u_cpu.rf_ram.memory\[121\]\[0\] _05935_ _05936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_204_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14406_ _00260_ net3 mod.u_cpu.rf_ram.memory\[484\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11618_ _02015_ _05218_ _05219_ _00702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_175_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15386_ _01161_ net3 mod.u_cpu.rf_ram.memory\[105\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_184_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12598_ _05890_ _01011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_102_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_156_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_204_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10223__A1 _04108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12236__I _03944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08967__A2 _03271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14337_ _00191_ net3 mod.u_cpu.rf_ram.memory\[51\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11549_ _05162_ mod.u_cpu.rf_ram.memory\[275\]\[1\] _05172_ _05174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_117_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14309__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10774__A2 _04225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14268_ _00122_ net3 mod.u_cpu.rf_ram.memory\[553\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_143_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08719__A2 mod.u_cpu.rf_ram.memory\[230\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13219_ _06317_ _06326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13712__A2 _06712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_252_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14199_ _03389_ mod.u_cpu.cpu.state.o_cnt\[2\] _07096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_174_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_174_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09545__I _03766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14459__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_98_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_239_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08760_ _02631_ _03059_ _03066_ _02363_ _03067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12523__I0 _05837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07711_ _01956_ _02011_ _02018_ _01989_ _02019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_39_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08691_ mod.u_cpu.rf_ram.memory\[200\]\[1\] mod.u_cpu.rf_ram.memory\[201\]\[1\] mod.u_cpu.rf_ram.memory\[202\]\[1\]
+ mod.u_cpu.rf_ram.memory\[203\]\[1\] _02349_ _02350_ _02998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_226_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_211_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07642_ mod.u_cpu.rf_ram.memory\[295\]\[0\] _01950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__13079__I1 _06221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09280__I _03495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_198_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07573_ _01663_ _01880_ _01881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_20_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09312_ _03557_ _03558_ _03560_ _03561_ _03562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10837__I0 _04682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_181_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08655__A1 _02124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12451__A2 _05788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_178_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_210_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09243_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[2\] _03503_ _03504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_181_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08750__S1 _02107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_221_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_210_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08407__A1 _02111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09174_ _03457_ _00016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12203__A2 _05611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_175_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08125_ _02405_ _02429_ _02432_ _02415_ _02433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__09080__A1 _03378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15234__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08056_ _02348_ _02351_ _02362_ _02363_ _02364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_190_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09907__A1 _03843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_192_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08499__C _02096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09383__A2 _03615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07233__I2 mod.u_cpu.rf_ram.memory\[458\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15384__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_130_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08958_ mod.u_cpu.cpu.decode.opcode\[2\] mod.u_cpu.cpu.decode.opcode\[0\] mod.u_cpu.cpu.decode.opcode\[1\]
+ _03263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XTAP_4615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_243_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_229_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11317__I1 mod.u_cpu.rf_ram.memory\[312\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3903 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07909_ _02216_ mod.u_cpu.rf_ram.memory\[208\]\[0\] _02217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_4659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3914 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3925 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08889_ mod.u_cpu.rf_ram.memory\[560\]\[1\] mod.u_cpu.rf_ram.memory\[561\]\[1\] mod.u_cpu.rf_ram.memory\[562\]\[1\]
+ mod.u_cpu.rf_ram.memory\[563\]\[1\] _02457_ _02473_ _03196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__07146__A1 _01452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_217_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_245_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_217_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3936 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3947 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10920_ _04743_ _00480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_99_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_217_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_205_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3958 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_16_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3969 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_186_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10851_ _04694_ _04695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_38_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11225__I _04951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_72_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08646__A1 _01670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_13570_ mod.u_arbiter.i_wb_cpu_dbus_adr\[18\] mod.u_arbiter.i_wb_cpu_dbus_adr\[19\]
+ _06604_ _06605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_201_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10782_ _04637_ mod.u_cpu.rf_ram.memory\[396\]\[0\] _04649_ _04650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_213_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_188_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_212_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_12521_ _05827_ mod.u_cpu.rf_ram.memory\[166\]\[0\] _05839_ _05840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XPHY_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__10453__A1 _04251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_234_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_125_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_197_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_240_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15240_ _01093_ net3 mod.u_cpu.rf_ram_if.rreq_r vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_12452_ _03394_ _05790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_185_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11253__I0 _04952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11403_ _04792_ _05058_ _05075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_172_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12056__I _05309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_184_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_15171_ _01024_ net3 mod.u_cpu.rf_ram.memory\[14\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_126_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12383_ _05741_ _00945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_158_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11953__A1 _05452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_193_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14122_ _03842_ _05631_ _07047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_126_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11334_ _04960_ _05028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_126_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_193_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14601__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09749__I1 _03929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14053_ mod.u_arbiter.i_wb_cpu_rdt\[26\] _06998_ _06993_ mod.u_arbiter.i_wb_cpu_dbus_dat\[26\]
+ _07002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_238_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11265_ _04980_ _00588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_106_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13004_ _01453_ _06172_ _03370_ _06173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_10216_ _04262_ _04263_ _04264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_106_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11196_ _04916_ mod.u_cpu.rf_ram.memory\[331\]\[1\] _04931_ _04933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_122_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13816__S _03510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10304__I _04248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10147_ _04068_ _04173_ _04213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_94_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14751__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_208_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14955_ _00809_ net3 mod.u_cpu.rf_ram.memory\[539\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_134_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_212_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10078_ _04142_ _04164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_208_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13906_ _06065_ _06490_ _06888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_36_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_14886_ _00740_ net3 mod.u_cpu.rf_ram.memory\[240\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08885__A1 _02500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_208_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_262_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13837_ _06340_ _06832_ _06833_ _01307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__15107__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_204_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_204_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13768_ _03674_ _06769_ _06770_ _06411_ _01301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_204_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13630__A1 _06485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12433__A2 _05774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_250_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_231_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_204_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08732__S1 _01525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12719_ _05970_ _01052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_15507_ _01278_ net3 mod.u_arbiter.i_wb_cpu_dbus_adr\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_203_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13699_ _03364_ _06704_ _06707_ _06708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__15257__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15438_ _01213_ net3 mod.u_cpu.rf_ram.memory\[139\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_248_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08444__I _01919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12197__A1 _05588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15369_ _01144_ net3 mod.u_cpu.rf_ram.memory\[108\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__13933__A2 mod.u_cpu.cpu.bufreg.lsb\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_184_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__14281__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09930_ _04002_ _04062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13697__A1 _06694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09861_ _04013_ _04014_ _04015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08812_ mod.u_cpu.rf_ram.memory\[12\]\[1\] mod.u_cpu.rf_ram.memory\[13\]\[1\] mod.u_cpu.rf_ram.memory\[14\]\[1\]
+ mod.u_cpu.rf_ram.memory\[15\]\[1\] _02266_ _02388_ _03119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_258_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10214__I _03950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09792_ _03963_ _00132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08743_ _02992_ _03011_ _03049_ _02148_ _03050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_113_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14110__A2 _05397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_227_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_213_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07679__A2 mod.u_cpu.rf_ram.memory\[278\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08674_ _02479_ mod.u_cpu.rf_ram.memory\[212\]\[1\] _02980_ _02981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_254_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_183_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07625_ mod.u_cpu.rf_ram.memory\[304\]\[0\] mod.u_cpu.rf_ram.memory\[305\]\[0\] mod.u_cpu.rf_ram.memory\[306\]\[0\]
+ mod.u_cpu.rf_ram.memory\[307\]\[0\] _01802_ _01932_ _01933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_199_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08628__A1 _02090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07556_ _01671_ _01864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__13621__A1 _06249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10884__I _04496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08723__S1 _01732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07487_ _01728_ mod.u_cpu.rf_ram.memory\[436\]\[0\] _01794_ _01795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_210_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09226_ _03488_ _03489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_107_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14177__A2 _03933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14624__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09157_ mod.u_arbiter.i_wb_cpu_rdt\[8\] _03436_ _03447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_213_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08108_ _02405_ _02409_ _02414_ _02415_ _02416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_163_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08800__A1 _03001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09088_ mod.u_cpu.cpu.state.o_cnt_r\[3\] _03389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_257_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08039_ _01630_ _02347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_135_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13688__A1 _06494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14774__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09185__I _03451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12735__I0 _05966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11050_ _04833_ _00520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09356__A2 _03586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09600__I0 _03800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_235_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07367__A1 _01670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_118_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10001_ _02529_ _04109_ _04110_ _00194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_5124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_130_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_114_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09913__I _04050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_218_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07861__C _02168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_184_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_3700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_218_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_4456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14740_ _00594_ net3 mod.u_cpu.rf_ram.memory\[317\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11952_ _03795_ _05452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_4489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08867__A1 _02461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_233_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_205_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13860__A1 _06465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10903_ _04731_ _00475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_244_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14671_ _00525_ net3 mod.u_cpu.rf_ram.memory\[352\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11883_ _05385_ mod.u_cpu.rf_ram.memory\[227\]\[0\] _05402_ _05403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_3799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_233_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_205_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13622_ _01935_ _06636_ _06637_ _01288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_73_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10834_ _04277_ _04669_ _04684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_260_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__12415__A2 _04228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_220_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_232_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_213_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11474__I0 _05108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13553_ _06595_ _01261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_242_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_198_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09292__A1 _03535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10765_ _04621_ _04637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_185_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_157_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12504_ _05827_ mod.u_cpu.rf_ram.memory\[16\]\[0\] _05828_ _05829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_157_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14168__A2 _06166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13484_ _03605_ _06545_ _06546_ _03610_ _06549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_40_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10696_ _04584_ mod.u_cpu.rf_ram.memory\[410\]\[0\] _04591_ _04592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__11226__I0 _04952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15223_ _01076_ net3 mod.u_cpu.rf_ram.memory\[131\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_172_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13915__A2 _06413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12435_ mod.u_cpu.rf_ram.memory\[173\]\[1\] _05765_ _05774_ _05776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_12_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_185_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11926__A1 _04994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11777__I1 mod.u_cpu.rf_ram.memory\[236\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15154_ _01007_ net3 mod.u_cpu.rf_ram.memory\[157\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12366_ _05730_ _00939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_154_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14105_ _03836_ _05720_ _07036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11317_ _05007_ mod.u_cpu.rf_ram.memory\[312\]\[0\] _05016_ _05017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_126_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15085_ _00939_ net3 mod.u_cpu.rf_ram.memory\[180\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_99_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12297_ _05139_ _05668_ _05683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08213__B _02520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11529__I1 mod.u_cpu.rf_ram.memory\[278\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07608__I _01581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14036_ _06914_ _06989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_11248_ _04968_ _00583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_136_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09028__C _03331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10201__I1 mod.u_cpu.rf_ram.memory\[48\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11179_ _04921_ _00561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_132_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08867__C _02578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_209_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_209_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_212_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_264_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_14938_ _00792_ net3 mod.u_cpu.rf_ram.memory\[223\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08858__A1 _01475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_236_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13851__A1 _06451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07343__I _01528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4990 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11701__I1 mod.u_cpu.rf_ram.memory\[252\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10665__A1 _03991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_263_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14869_ _00723_ net3 mod.u_cpu.rf_ram.memory\[255\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_1_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07410_ _01703_ _01708_ _01715_ _01717_ _01718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_23_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08375__S _02585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08390_ _02272_ _02696_ _02697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_95_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_177_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14647__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07341_ _01647_ _01648_ _01649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09283__A1 _03528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_189_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10968__A2 _04759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14159__A2 _03270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07272_ _01578_ _01579_ _01580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_176_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_223_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09011_ mod.u_cpu.cpu.bufreg.lsb\[0\] _03292_ _03316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_192_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_178_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11217__I0 _04938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13906__A2 _06490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09035__A1 _03338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_191_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__14797__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07946__C _01766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_258_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07597__A1 _01875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10440__I1 mod.u_cpu.rf_ram.memory\[452\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07518__I _01825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09934__S _04063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09913_ _04050_ _04051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_63_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12342__A1 _05494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09844_ _03752_ _04003_ _04004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_58_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_259_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08777__C _01916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09775_ _03950_ _03951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_3007 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14095__A1 _03804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3018 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08726_ _02161_ mod.u_cpu.rf_ram.memory\[244\]\[1\] _03032_ _03033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_3029 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08849__A1 _03001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08349__I _01841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_170_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15422__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13842__A1 mod.u_cpu.cpu.immdec.imm24_20\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_227_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07253__I _01560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_255_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_226_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_215_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08657_ _02104_ _02963_ _02964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_15_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_199_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_187_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_215_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_230_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07608_ _01581_ _01916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_1638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_242_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_202_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08588_ mod.u_cpu.rf_ram.memory\[269\]\[1\] _02895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_183_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_263_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_214_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07539_ _01836_ _01846_ _01485_ _01847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__15572__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11503__I _04959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_210_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10550_ _04481_ mod.u_cpu.rf_ram.memory\[434\]\[1\] _04491_ _04493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_195_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_224_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11208__I0 _04936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09209_ _03477_ _00033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_127_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_167_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10481_ _04436_ _04447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_120_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12220_ _05629_ _05630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_68_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07588__A1 _01893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11384__A2 _04779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12151_ _05583_ mod.u_cpu.rf_ram.memory\[207\]\[1\] _05580_ _05584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_2_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_194_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08880__S0 _02494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_190_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08033__B _02321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11102_ _04868_ _04869_ _04870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_155_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12082_ _05537_ _00848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_96_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12333__A1 _03879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08968__B mod.u_cpu.cpu.immdec.imm24_20\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11033_ _03959_ _04821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_110_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08632__S0 _02092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_249_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07591__C _01867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_218_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12984_ _06157_ _01130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_4286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_218_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14723_ _00577_ net3 mod.u_cpu.rf_ram.memory\[326\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11935_ _05440_ _00798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_27_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_245_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_233_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_233_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11614__S _05215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14654_ _00508_ net3 mod.u_cpu.rf_ram.memory\[360\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_60_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11866_ _05383_ mod.u_cpu.rf_ram.memory\[70\]\[1\] _05389_ _05391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_150_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_261_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_162_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2895 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13605_ _03362_ _03354_ _06624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_10817_ _04262_ _04669_ _04673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_159_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14585_ _00439_ net3 mod.u_cpu.rf_ram.memory\[395\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_198_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13061__A2 _06209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11797_ _03931_ _05343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_9_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_242_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13536_ mod.u_arbiter.i_wb_cpu_dbus_adr\[3\] mod.u_arbiter.i_wb_cpu_dbus_adr\[4\]
+ _06584_ _06586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07815__A2 _02108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10748_ _04626_ mod.u_cpu.rf_ram.memory\[402\]\[1\] _04624_ _04627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_159_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13467_ _06537_ _06538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_127_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10679_ _04307_ _04570_ _04581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_15206_ _01059_ net3 mod.u_cpu.rf_ram.memory\[209\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_173_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12418_ _05229_ _05765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09568__A2 _03747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13398_ _06285_ _06492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11375__A2 _05055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15137_ _00990_ net3 mod.u_cpu.rf_ram.memory\[429\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_154_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12349_ _05718_ _00934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_99_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07338__I _01645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_141_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15068_ _00922_ net3 mod.u_cpu.rf_ram.memory\[185\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_142_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12175__I1 mod.u_cpu.rf_ram.memory\[76\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08878__B _03184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_253_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14019_ mod.u_arbiter.i_wb_cpu_rdt\[17\] _06976_ _06971_ mod.u_arbiter.i_wb_cpu_dbus_dat\[17\]
+ _06977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_07890_ _02197_ _02198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08623__S0 _01925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15445__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_255_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14077__A1 _03910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13124__I0 _06237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09560_ _03749_ _03779_ _03780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_209_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_237_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08511_ mod.u_cpu.rf_ram.memory\[350\]\[1\] mod.u_cpu.rf_ram.memory\[351\]\[1\] _01664_
+ _02818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_110_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_224_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_209_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_208_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11686__I0 _05250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_184_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09491_ mod.u_cpu.rf_ram_if.wen1_r mod.u_cpu.rf_ram_if.wen0_r _01418_ _03717_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_36_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07503__A1 _01773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15595__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13803__I _06424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08442_ mod.u_cpu.rf_ram.memory\[392\]\[1\] mod.u_cpu.rf_ram.memory\[393\]\[1\] mod.u_cpu.rf_ram.memory\[394\]\[1\]
+ mod.u_cpu.rf_ram.memory\[395\]\[1\] _02020_ _02748_ _02749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_224_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_208_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07801__I _01701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11438__I0 _05096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08373_ _01591_ _02653_ _02679_ _02680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_260_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_189_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_221_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07324_ _01631_ _01632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_220_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07806__A2 mod.u_cpu.rf_ram.memory\[172\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_192_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07255_ _01561_ _01562_ _01563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_176_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_149_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07186_ mod.u_cpu.raddr\[0\] _01494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_105_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12563__A1 _05417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_258_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_219_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07248__I _01539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09664__S _03860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08909__I2 mod.u_cpu.rf_ram.memory\[522\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_150_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08614__S0 _02059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09827_ _03989_ _00141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10877__A1 _04611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14812__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08300__C _02606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_228_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09758_ _03936_ mod.u_cpu.rf_ram.memory\[552\]\[1\] _03934_ _03937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_73_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_251_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_261_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_215_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08709_ _02594_ _03012_ _03015_ _02764_ _03016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XTAP_2114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_104_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_227_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09689_ _03862_ mod.u_cpu.rf_ram.memory\[55\]\[1\] _03880_ _03882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09495__A1 _03374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11720_ _05037_ _05284_ _05290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_230_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_243_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_203_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14962__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13418__I1 mod.u_cpu.rf_ram.memory\[339\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_230_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11429__I0 _05087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11651_ _05234_ mod.u_cpu.rf_ram.memory\[24\]\[1\] _05240_ _05242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_168_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_147_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_230_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10602_ _03892_ _04225_ _04528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_14370_ _00224_ net3 mod.u_cpu.rf_ram.memory\[502\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11582_ _05110_ _03797_ _05196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_70_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_196_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13321_ _06417_ _06418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_156_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15318__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_182_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10533_ _04481_ mod.u_cpu.rf_ram.memory\[437\]\[1\] _04479_ _04482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_210_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_182_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09638__I _03841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12929__I0 _06107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13252_ _04984_ _06344_ _06352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10464_ _04434_ _00333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_237_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12203_ _05343_ _05611_ _05619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_164_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13751__B1 _06326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10404__I1 mod.u_cpu.rf_ram.memory\[458\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13183_ _03500_ mod.u_arbiter.i_wb_cpu_rdt\[5\] _06290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_159_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10395_ _03727_ _03807_ _04389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_163_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15468__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14342__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12134_ _05334_ _05543_ _05572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_150_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13096__S _06231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07981__A1 _02135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12065_ _02395_ _05525_ _05526_ _00842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_123_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_237_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11016_ _04803_ mod.u_cpu.rf_ram.memory\[35\]\[0\] _04809_ _04810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_49_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14492__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08081__S1 _02388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11408__I _03712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_253_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4050 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_168_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4061 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13806__A1 _06735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4072 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_161_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_219_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13806__B2 _06332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_206_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4083 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4094 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09486__A1 _03702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08289__A2 _02595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12967_ _03338_ _03375_ _06143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_3371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_206_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11293__A1 _04859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14706_ _00560_ net3 mod.u_cpu.rf_ram.memory\[334\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11918_ _03750_ _05428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_3393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_209_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10340__I0 _04345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12898_ _06072_ _06088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_2670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_220_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_209_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_206_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07621__I _01686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10891__I1 _04661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11849_ _05366_ mod.u_cpu.rf_ram.memory\[149\]\[0\] _05378_ _05379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_14637_ _00491_ net3 mod.u_cpu.rf_ram.memory\[36\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_221_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_221_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_207_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1980 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1991 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_158_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09749__S _03926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12093__I0 _05539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14568_ _00422_ net3 mod.u_cpu.rf_ram.memory\[403\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_18_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08836__I1 mod.u_cpu.rf_ram.memory\[49\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_174_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_118_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10643__I1 _04532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13519_ _06568_ _03691_ _06572_ _06573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_14499_ _00353_ net3 mod.u_cpu.rf_ram.memory\[438\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_88_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09548__I _03769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_256_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08452__I _01615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_161_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_177_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_216_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08991_ _03260_ _03294_ _03295_ _03296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_130_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14835__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07972__A1 _02148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07942_ mod.u_cpu.rf_ram.memory\[239\]\[0\] _02250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_141_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_229_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10859__A1 mod.u_cpu.cpu.immdec.imm11_7\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07873_ mod.u_cpu.rf_ram.memory\[207\]\[0\] _02181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__07724__A1 _01997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_214_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09612_ _03821_ _03822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_96_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_256_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_243_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__14985__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09543_ _03765_ _00081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_71_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09477__A1 _01439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__13533__I _06583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12320__I1 mod.u_cpu.rf_ram.memory\[189\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_221_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_212_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09474_ _01418_ _01645_ _03700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_225_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_169_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_212_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_196_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08425_ _02687_ _02723_ _02731_ _01678_ _02732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__09229__A1 _03410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_180_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13025__A2 _06080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_212_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08356_ _02631_ _02662_ _01618_ _02663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_20_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07307_ _01614_ _01615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08287_ _02030_ _02594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_137_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_192_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_192_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14365__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07238_ mod.u_cpu.rf_ram.memory\[463\]\[0\] _01546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_180_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15610__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12536__A1 _05226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08204__A2 mod.u_cpu.rf_ram.memory\[564\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07169_ _01477_ _00007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08835__S0 _02151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09952__A2 _04077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10180_ _03910_ _04238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_133_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07963__A1 _02244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10333__S _04342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12839__A2 _06048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_219_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11228__I _03924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13870_ _06861_ _06862_ _06863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_47_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12821_ _06037_ _01087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_264_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_27_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_216_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_167_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12752_ _05991_ _01064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_15540_ _01311_ net3 mod.u_cpu.cpu.immdec.imm24_20\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_199_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_231_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_202_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11703_ _05271_ mod.u_cpu.rf_ram.memory\[252\]\[1\] _05276_ _05278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_203_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15140__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15471_ _01245_ net3 mod.u_cpu.cpu.ctrl.o_ibus_adr\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_203_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12683_ _05946_ _01040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14422_ _00276_ net3 mod.u_cpu.rf_ram.memory\[476\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11634_ mod.u_cpu.rf_ram.memory\[261\]\[1\] _05230_ _05227_ _05231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__14708__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_196_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13972__B1 _06919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14353_ _00207_ net3 mod.u_cpu.rf_ram.memory\[511\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11565_ _05180_ mod.u_cpu.rf_ram.memory\[272\]\[0\] _05184_ _05185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__11822__I0 _05342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_183_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08443__A2 _02749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13304_ _06118_ _06300_ _06402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__15290__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10516_ _04471_ _00348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_14284_ _00138_ net3 mod.u_cpu.rf_ram.memory\[545\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_109_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11496_ _05138_ _00661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_171_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12527__A1 _05843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14858__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13235_ _03751_ _06193_ _06341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_108_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10447_ _04347_ _04423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_136_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_13166_ _06275_ _01194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_10378_ _04376_ _00305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_112_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07954__A1 _02180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12117_ _05559_ mod.u_cpu.rf_ram.memory\[210\]\[0\] _05560_ _05561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_2_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10243__S _04282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13097_ _06233_ _01167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07616__I _01634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_215_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12048_ _05514_ _00837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_78_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07706__A1 _01998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13781__C _06432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_225_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_168_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14238__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_207_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13999_ _06960_ _06961_ _01341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_94_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_222_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_207_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10313__I0 _04326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_234_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07351__I mod.u_cpu.raddr\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_206_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07565__S0 _01843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_221_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14204__A1 _06153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13007__A2 _06080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_181_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08210_ _02291_ _02518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__14388__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12066__I0 _05518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_222_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09190_ mod.u_arbiter.i_wb_cpu_rdt\[21\] mod.u_arbiter.i_wb_cpu_dbus_dat\[18\] _03464_
+ _03467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_194_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15633__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_147_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08141_ _02124_ _02449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_53_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13302__B _06381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11813__I0 _05350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08434__A2 _02733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08072_ _01485_ _02380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_31_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08985__A3 mod.u_cpu.cpu.state.o_cnt_r\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08198__A1 _02449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07945__A1 _02249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_248_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08974_ mod.u_cpu.cpu.bufreg.lsb\[0\] _03279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__15013__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07925_ mod.u_cpu.rf_ram.memory\[224\]\[0\] mod.u_cpu.rf_ram.memory\[225\]\[0\] mod.u_cpu.rf_ram.memory\[226\]\[0\]
+ mod.u_cpu.rf_ram.memory\[227\]\[0\] _02151_ _02172_ _02233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_4808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_151_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_130_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_229_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07856_ _01820_ _02164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_57_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09741__I _03696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_217_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07173__A2 _01479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15163__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07787_ _02090_ _02094_ _02095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_83_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09526_ _03745_ _03749_ _03750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__07261__I _01568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_149_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09170__I0 mod.u_arbiter.i_wb_cpu_rdt\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_266_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09457_ _03356_ _03680_ _03682_ _03684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_101_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_200_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__11009__A1 _04804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08408_ _02462_ mod.u_cpu.rf_ram.memory\[444\]\[1\] _02714_ _02715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_197_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09388_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[24\] mod.u_cpu.cpu.ctrl.o_ibus_adr\[23\] mod.u_cpu.cpu.ctrl.o_ibus_adr\[22\]
+ _03606_ _03626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_177_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_200_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08339_ _02421_ _02645_ _02646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_138_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12607__I _04024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11511__I _05124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_193_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11350_ _05028_ mod.u_cpu.rf_ram.memory\[307\]\[0\] _05039_ _05040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_197_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11280__I1 mod.u_cpu.rf_ram.memory\[318\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12509__A1 _05343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08025__C _01717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10301_ _04324_ _00280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_11281_ _04992_ _00592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_180_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_152_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13020_ _06183_ _01140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_106_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_238_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10232_ _04267_ mod.u_cpu.rf_ram.memory\[484\]\[1\] _04273_ _04275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09925__A2 _03843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10163_ _04223_ _04224_ _04225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__07436__I _01743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_266_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14971_ _00825_ net3 mod.u_cpu.rf_ram.memory\[57\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10094_ _01597_ _04174_ _04175_ _00222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_130_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08036__S1 _01638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15506__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13922_ _06166_ _06649_ _06900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_43_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_207_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07164__A2 mod.u_cpu.cpu.immdec.imm19_12_20\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_262_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13853_ mod.u_cpu.cpu.immdec.imm24_20\[1\] _06836_ _06837_ mod.u_cpu.cpu.immdec.imm24_20\[2\]
+ _06848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_12804_ _06019_ mod.u_cpu.rf_ram.memory\[128\]\[1\] _06024_ _06026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_250_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14530__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07171__I mod.u_cpu.cpu.immdec.imm19_12_20\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13784_ _06065_ _06783_ _06785_ _06786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_10996_ _03761_ _04795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_203_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_204_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15523_ _01294_ net3 mod.u_cpu.cpu.immdec.imm19_12_20\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_167_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09456__A4 _03682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12735_ _05966_ mod.u_cpu.rf_ram.memory\[136\]\[1\] _05979_ _05981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09861__A1 _04013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_241_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_163_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_231_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_176_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15454_ _01228_ net3 mod.u_cpu.cpu.ctrl.o_ibus_adr\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12666_ _05896_ _05721_ _05935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_231_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_129_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_204_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12748__A1 _05395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11617_ _05133_ _05218_ _05219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__14680__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14405_ _00259_ net3 mod.u_cpu.rf_ram.memory\[485\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_204_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15385_ _01160_ net3 mod.u_cpu.rf_ram.memory\[105\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_30_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12597_ _05887_ mod.u_cpu.rf_ram.memory\[155\]\[0\] _05889_ _05890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_50_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11420__A1 _05022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10223__A2 _04228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11548_ _05173_ _00678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_184_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14336_ _00190_ net3 mod.u_cpu.rf_ram.memory\[51\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_183_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_239_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14267_ _00121_ net3 mod.u_cpu.rf_ram.memory\[554\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_143_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11479_ _05114_ mod.u_cpu.rf_ram.memory\[286\]\[0\] _05126_ _05127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_171_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15036__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13173__A1 mod.u_cpu.cpu.bufreg.i_sh_signed vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13218_ _06307_ _06315_ _06319_ _06324_ _06325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_174_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14198_ _07076_ _03320_ _01406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__07927__A1 _02157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_258_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12920__A1 _05888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_170_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13149_ _06265_ _01187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_3_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12771__I1 _05971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10782__I0 _04637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_174_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_257_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15186__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07710_ _01961_ _02014_ _02017_ _02005_ _02018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_254_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_266_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08690_ _02578_ _02993_ _02996_ _02660_ _02997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_250_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09561__I _03780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08352__A1 _02656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07786__S0 _02092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07641_ _01758_ _01949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_66_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_253_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07572_ mod.u_cpu.rf_ram.memory\[375\]\[0\] _01880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07538__S0 _01832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09311_ _03486_ _03561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_22_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08655__A2 _02954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09242_ _03502_ _03503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_142_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_194_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09173_ _03456_ mod.u_arbiter.i_wb_cpu_dbus_dat\[11\] _03452_ _03457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08407__A2 _02713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08124_ _02410_ mod.u_cpu.rf_ram.memory\[38\]\[0\] _02431_ _01828_ _02432_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_175_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_190_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08055_ _01586_ _02363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_134_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09368__B1 _03401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13164__A1 _05515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09907__A2 _04038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14403__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15529__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_142_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_249_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09672__S _03867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08591__A1 _02759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08957_ mod.u_cpu.cpu.decode.co_ebreak _01423_ _03262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_217_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11478__A1 _04852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07908_ _01681_ _02216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_4649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3904 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08888_ _02449_ _03187_ _03194_ _02505_ _03195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__10525__I0 _04469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14553__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3915 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_99_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09471__I _03696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3926 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07146__A2 _01454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08343__A1 _02638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_244_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3937 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3948 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07839_ _02103_ _02146_ _01475_ _02147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_99_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3959 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_72_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12278__I0 _05660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10850_ _04620_ _04694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_232_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_232_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09509_ _03733_ _03734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10781_ _04233_ _04648_ _04649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_227_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12520_ _05355_ _05831_ _05839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_80_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_201_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__10453__A2 _03905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_198_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__07859__C _02166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_200_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_185_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_205_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_185_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12451_ _03700_ _05788_ _05789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_184_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12337__I _05709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10058__S _04149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_227_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15059__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11402_ _05074_ _00631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_166_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_15170_ _01023_ net3 mod.u_cpu.rf_ram.memory\[14\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_138_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12382_ _05729_ mod.u_cpu.rf_ram.memory\[178\]\[1\] _05739_ _05741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_181_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14121_ _07046_ _01378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_11333_ _05027_ _00609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11953__A2 _05423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_181_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14052_ mod.u_arbiter.i_wb_cpu_dbus_dat\[27\] _07000_ _07001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11264_ _04978_ mod.u_cpu.rf_ram.memory\[320\]\[0\] _04979_ _04980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_125_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07909__A1 _02216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13003_ _01435_ _01420_ _01424_ _06172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_234_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10215_ _04136_ _04263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_11195_ _04932_ _00566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08582__A1 _02027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07166__I _01474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_239_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10146_ _04212_ _00237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_121_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_43_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14954_ _00808_ net3 mod.u_cpu.rf_ram.memory\[539\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10077_ _04025_ _04163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_48_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__08334__A1 _02638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_263_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_13905_ _06481_ _06660_ _06887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_78_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14885_ _00739_ net3 mod.u_cpu.rf_ram.memory\[241\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_78_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_235_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_223_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13836_ mod.u_cpu.cpu.immdec.imm30_25\[5\] _06774_ _06833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_251_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_3 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_245_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13767_ _06764_ _03391_ _06416_ _06770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_10979_ _04783_ _00499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_189_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13630__A2 _06284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_189_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15506_ _01277_ net3 mod.u_arbiter.i_wb_cpu_dbus_adr\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12718_ _05966_ mod.u_cpu.rf_ram.memory\[138\]\[1\] _05968_ _05970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_91_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_231_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13698_ _06421_ _06706_ _06707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_31_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12247__I _03967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15437_ _01212_ net3 mod.u_cpu.rf_ram.memory\[91\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_129_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12649_ _05924_ _01028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_102_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12197__A2 _05594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13394__A1 _06485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_200_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_156_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15368_ _01143_ net3 mod.u_cpu.rf_ram.memory\[84\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__14426__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14319_ _00173_ net3 mod.u_cpu.rf_ram.memory\[528\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_183_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15299_ _00059_ net4 mod.u_scanchain_local.module_data_in\[56\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_116_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_264_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_252_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__13078__I _03734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13697__A2 _06431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_259_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09860_ _03836_ _04014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14576__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_217_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08573__A1 _01949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08811_ mod.u_cpu.rf_ram.memory\[0\]\[1\] mod.u_cpu.rf_ram.memory\[1\]\[1\] mod.u_cpu.rf_ram.memory\[2\]\[1\]
+ mod.u_cpu.rf_ram.memory\[3\]\[1\] _02211_ _02386_ _03118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09791_ _03958_ mod.u_cpu.rf_ram.memory\[548\]\[0\] _03962_ _03963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_100_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10380__A1 _03721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08742_ _01848_ _03029_ _03048_ _03049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_226_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08673_ _02202_ _02979_ _02980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_113_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08876__A2 mod.u_cpu.rf_ram.memory\[558\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_227_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_214_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07624_ _01827_ _01932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_187_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_214_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12866__B _06046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07555_ _01862_ _01863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_241_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08628__A2 _02934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_222_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15201__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_224_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12680__I0 _05934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07486_ _01774_ _01793_ _01794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07679__C _01952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_194_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13909__B1 _06443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09225_ _03487_ _03488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_167_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_194_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13385__A1 _06397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09156_ mod.u_arbiter.i_wb_cpu_dbus_dat\[5\] _03446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_135_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08107_ _01765_ _02415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__15351__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09087_ mod.u_cpu.cpu.state.o_cnt_r\[0\] _03388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_163_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10994__I0 _04774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_194_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_190_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14919__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09466__I _03692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14185__I0 _07081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_174_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08370__I _01886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08038_ _02339_ _02341_ _02343_ _02345_ _02346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__13688__A2 _06644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_235_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08564__A1 _01961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07367__A2 _01674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10000_ _03899_ _04109_ _04110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_49_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_130_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09989_ _04091_ mod.u_cpu.rf_ram.memory\[51\]\[1\] _04100_ _04102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_114_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_218_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13716__I _05784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_123_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08316__A1 _02566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_188_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07714__I _01704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_218_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_4468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11951_ _05451_ _00803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10123__A1 _04196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_218_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_217_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11236__I _04959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13860__A2 _06744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_123_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10902_ _04720_ mod.u_cpu.rf_ram.memory\[377\]\[1\] _04729_ _04731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_11882_ _04965_ _05401_ _05402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_3778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14670_ _00524_ net3 mod.u_cpu.rf_ram.memory\[352\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_264_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_13621_ _06249_ _06636_ _06637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_60_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10833_ _04683_ _00453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_53_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_242_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_41_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11623__A1 _04812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_186_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08545__I _01886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10764_ _04636_ _00431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_13552_ mod.u_arbiter.i_wb_cpu_dbus_adr\[10\] mod.u_arbiter.i_wb_cpu_dbus_adr\[11\]
+ _06594_ _06595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12671__I0 _05938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_213_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14449__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_197_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12503_ _05563_ _03873_ _05828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_125_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_13483_ _06548_ _01238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_201_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_200_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10695_ _04322_ _04575_ _04591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_139_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15222_ _01075_ net3 mod.u_cpu.rf_ram.memory\[131\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12434_ _02112_ _05774_ _05775_ _00962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11226__I1 mod.u_cpu.rf_ram.memory\[326\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12423__I0 _05753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_194_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13099__S _06234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_201_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12365_ _05729_ mod.u_cpu.rf_ram.memory\[180\]\[1\] _05727_ _05730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_15153_ _01006_ net3 mod.u_cpu.rf_ram.memory\[158\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_201_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14599__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09376__I _03614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11316_ _04732_ _05011_ _05016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_153_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14104_ _07035_ _01372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_153_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15084_ _00938_ net3 mod.u_cpu.rf_ram.memory\[180\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_181_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12296_ _05682_ _00917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_180_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14035_ _06986_ _06988_ _01350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_4_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11247_ _04952_ mod.u_cpu.rf_ram.memory\[323\]\[1\] _04966_ _04968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_175_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08555__A1 _01981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11178_ _04916_ mod.u_cpu.rf_ram.memory\[334\]\[1\] _04919_ _04921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_80_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10362__A1 _04209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_209_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10129_ _03858_ _04201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_110_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07624__I _01827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08307__A1 _02566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_208_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14937_ _00791_ net3 mod.u_cpu.rf_ram.memory\[224\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10114__A1 _04189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_224_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08858__A2 _03141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4980 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_180_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4991 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13851__A2 _06672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_224_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10665__A2 _04570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15224__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14868_ _00722_ net3 mod.u_cpu.rf_ram.memory\[255\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_63_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_223_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_13819_ _06363_ _06465_ _06668_ _06779_ _06818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_189_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14799_ _00653_ net3 mod.u_cpu.rf_ram.memory\[288\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_91_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_211_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08166__S0 _02472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_250_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07340_ mod.u_cpu.rf_ram.memory\[495\]\[0\] _01648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_188_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_204_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07271_ mod.u_cpu.rf_ram.memory\[471\]\[0\] _01579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__15374__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_176_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09010_ _01428_ _03315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_148_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_191_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_145_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08794__A1 _02202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07597__A2 mod.u_cpu.rf_ram.memory\[356\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09912_ _03738_ _04050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_176_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10728__I0 _04608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08546__A1 _02196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12342__A2 _05703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09843_ _04002_ _04003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_99_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_112_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_258_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_219_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_230_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09774_ _03949_ _03950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_86_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14095__A2 _07014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3008 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3019 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_227_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08725_ _02197_ _03031_ _03032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_227_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11153__I0 _04896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13842__A2 _06836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_254_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11853__A1 _05239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08656_ _02105_ _02953_ _02962_ _02963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_2329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10900__I0 _04728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_265_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_265_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07607_ _01914_ _01915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_82_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08587_ mod.u_cpu.rf_ram.memory\[270\]\[1\] mod.u_cpu.rf_ram.memory\[271\]\[1\] _02106_
+ _02894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_41_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_228_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11605__A1 _05078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07538_ _01839_ _01840_ _01842_ _01845_ _01832_ _01833_ _01846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__08365__I _02026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12653__I0 _05923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07469_ _01728_ mod.u_cpu.rf_ram.memory\[428\]\[0\] _01776_ _01777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_183_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12816__S _06031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_249_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13358__A1 _06395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14741__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09208_ mod.u_arbiter.i_wb_cpu_rdt\[29\] mod.u_arbiter.i_wb_cpu_dbus_dat\[26\] _03474_
+ _03477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_127_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12405__I0 _05745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10480_ _04446_ _00337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_176_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_202_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09139_ mod.u_arbiter.i_wb_cpu_dbus_dat\[1\] _03433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_108_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_191_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07588__A2 mod.u_cpu.rf_ram.memory\[364\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08785__A1 _01696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12150_ _05549_ _05583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_191_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08880__S1 _02451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11101_ _04847_ _04869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_155_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14891__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12081_ _05521_ mod.u_cpu.rf_ram.memory\[212\]\[0\] _05536_ _05537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12551__S _05856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10719__I0 _04598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11032_ _04820_ _00515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12333__A2 _05703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10344__A1 _04352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11392__I0 _05046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13446__I _06510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08632__S1 _02098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_77_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_4221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15247__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07444__I _01645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12097__A1 _04965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12983_ mod.u_cpu.cpu.genblk3.csr.mstatus_mie mod.u_cpu.cpu.genblk3.csr.mstatus_mpie
+ _06143_ _06157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_4276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13833__A2 _06829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08984__B _01421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14722_ _00576_ net3 mod.u_cpu.rf_ram.memory\[326\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11934_ mod.u_cpu.rf_ram.memory\[169\]\[0\] _05437_ _05439_ _05440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_3564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14271__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_205_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__15397__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14653_ _00507_ net3 mod.u_cpu.rf_ram.memory\[361\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11865_ _05390_ _00778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_260_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__15313__D mod.u_scanchain_local.module_data_in\[69\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2896 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_232_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13604_ _06623_ _01284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13597__A1 _03659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10816_ _04672_ _00447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_11796_ _05310_ _05342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_14584_ _00438_ net3 mod.u_cpu.rf_ram.memory\[395\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_198_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08208__C _02515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13535_ _06585_ _01253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_10747_ _04578_ _04626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_201_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_127_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10678_ _04580_ _00401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_13466_ _06509_ _06537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09017__A2 mod.u_cpu.cpu.ctrl.i_iscomp vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_185_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_145_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15205_ _01058_ net3 mod.u_cpu.rf_ram.memory\[136\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12417_ _05764_ _00956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_127_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13397_ _06478_ _06479_ _06481_ _06491_ _01209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__10958__I0 _04756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08776__A1 _01863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15136_ _00989_ net3 mod.u_cpu.rf_ram.memory\[429\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_114_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_126_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12348_ _05713_ mod.u_cpu.rf_ram.memory\[181\]\[0\] _05717_ _05718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_173_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15067_ _00921_ net3 mod.u_cpu.rf_ram.memory\[186\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_99_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12279_ _05671_ _00911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_114_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08528__A1 _01977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09834__I _03995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14018_ _06963_ _06976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08878__C _01836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13356__I _06426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08623__S1 _02071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_256_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__14077__A2 _04996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07354__I _01661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09770__S _03943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_209_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_209_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14614__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_255_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_236_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08510_ _02664_ _02807_ _02816_ _02817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_48_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09490_ _03664_ _03715_ _03716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_64_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_252_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08700__A1 _01573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07503__A2 _01805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08441_ _01762_ _02748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_1_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_247_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_224_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14764__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08372_ _02661_ _02663_ _02664_ _02678_ _02679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_251_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_225_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07323_ _01630_ _01631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07267__A1 _01573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12260__A1 _05657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_177_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_192_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07254_ mod.u_cpu.rf_ram.memory\[479\]\[0\] _01562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_164_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07957__C _02168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_191_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07185_ _01492_ _01493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_121_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_219_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07529__I _01510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08767__A1 _02303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13760__A1 mod.u_cpu.cpu.immdec.imm31 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12563__A2 _05757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07973__B _01481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_259_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08614__S1 _01723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_232_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_189_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09826_ _03964_ mod.u_cpu.rf_ram.memory\[544\]\[1\] _03987_ _03989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_24_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07264__I _01504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_228_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_150_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14294__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09757_ _03889_ _03936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_215_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_215_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_255_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11826__A1 _04294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08708_ _02209_ _03013_ _03014_ _02633_ _03015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XTAP_2115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_215_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09688_ _03881_ _00110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_15_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08639_ mod.u_cpu.rf_ram.memory\[173\]\[1\] _02946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_242_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11650_ _05241_ _00712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_214_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_199_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11429__I1 mod.u_cpu.rf_ram.memory\[294\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_120_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_168_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10601_ _03713_ _04527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_35_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11581_ _05195_ _00689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_70_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08845__I2 mod.u_cpu.rf_ram.memory\[42\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_195_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13320_ _06313_ _06417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_168_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10532_ _04429_ _04481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_161_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__12929__I1 mod.u_cpu.rf_ram.memory\[369\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10463_ _04430_ mod.u_cpu.rf_ram.memory\[448\]\[1\] _04432_ _04434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_109_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13251_ _06204_ _06351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_202_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_182_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08758__A1 _02204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07439__I _01746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12202_ _05618_ _00887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13751__B2 _06281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13182_ _06288_ _06289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_136_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10394_ _04388_ _00309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_191_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10565__A1 _04369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12133_ _05571_ _00865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_151_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_150_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12064_ _05488_ _05525_ _05526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_150_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14637__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13176__I _06282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11015_ _04808_ _03969_ _04809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_104_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_238_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08930__A1 _02509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4040 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_213_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4051 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_237_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4062 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_218_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4073 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_218_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4084 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4095 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14787__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12966_ _01425_ _06142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_234_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09486__A2 _03711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_248_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14705_ _00559_ net3 mod.u_cpu.rf_ram.memory\[335\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11917_ _05427_ _00793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07497__A1 _01517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10340__I1 mod.u_cpu.rf_ram.memory\[468\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12897_ _06087_ _01113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_261_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_178_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_233_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_221_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14636_ _00490_ net3 mod.u_cpu.rf_ram.memory\[36\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_53_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11848_ _04014_ _05374_ _05378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_127_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1970 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1981 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_202_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1992 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12242__A1 _05367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_207_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13290__I0 mod.u_arbiter.i_wb_cpu_rdt\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14567_ _00421_ net3 mod.u_cpu.rf_ram.memory\[404\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11779_ _04930_ _05301_ _05331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_220_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13518_ _03685_ _03690_ _06572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_140_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14498_ _00352_ net3 mod.u_cpu.rf_ram.memory\[438\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_158_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13449_ _06527_ _01225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__13042__I0 _06186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08749__A1 _02611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15412__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13287__S _06377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15119_ _00972_ net3 mod.u_cpu.rf_ram.memory\[449\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_47_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__10704__S _04595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08990_ _03278_ _03293_ _03267_ _03295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_86_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_253_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07941_ _01539_ _02249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_130_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__15562__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08401__C _01981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07872_ _01778_ _02180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_25_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08921__A1 _02528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09611_ _03818_ _03820_ _03821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_28_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09542_ _03764_ mod.u_cpu.rf_ram.memory\[574\]\[1\] _03759_ _03765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_110_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09477__A2 _01494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09721__I0 _03890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09473_ _03698_ _03699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12481__A1 _05657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_224_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_52_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_197_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08424_ _02611_ _02726_ _02729_ _02730_ _02731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_145_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_260_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_200_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08355_ mod.u_cpu.rf_ram.memory\[488\]\[1\] mod.u_cpu.rf_ram.memory\[489\]\[1\] mod.u_cpu.rf_ram.memory\[490\]\[1\]
+ mod.u_cpu.rf_ram.memory\[491\]\[1\] _02385_ _02633_ _02662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__08288__I0 mod.u_cpu.rf_ram.memory\[456\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_177_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07306_ _01523_ _01614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_149_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08988__A1 _03279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_220_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08286_ _02116_ _02593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_177_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07237_ _01516_ _01545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_192_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13033__I0 _06184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15092__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12536__A2 _05438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07168_ _01447_ _01459_ _01466_ _01476_ _01477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_118_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10547__A1 _04201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08835__S1 _02152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_160_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07963__A2 mod.u_cpu.rf_ram.memory\[252\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08311__C _01742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_232_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08912__A1 _02546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09809_ _03958_ mod.u_cpu.rf_ram.memory\[546\]\[0\] _03976_ _03977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09960__I0 _04071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_219_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12820_ _06035_ mod.u_cpu.rf_ram.memory\[126\]\[0\] _06036_ _06037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_43_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12751_ _05984_ mod.u_cpu.rf_ram.memory\[199\]\[1\] _05989_ _05991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_257_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_203_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_243_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11702_ _05277_ _00728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_163_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08771__S0 _01664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15470_ _01244_ net3 mod.u_cpu.cpu.ctrl.o_ibus_adr\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12682_ _05938_ mod.u_cpu.rf_ram.memory\[142\]\[1\] _05944_ _05946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_203_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_231_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14421_ _00275_ net3 mod.u_cpu.rf_ram.memory\[477\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12224__A1 _02330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11633_ _05229_ _05230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08279__I0 mod.u_cpu.rf_ram.memory\[462\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_243_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_202_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09649__I _03850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10086__I0 _04162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15435__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14352_ _00206_ net3 mod.u_cpu.rf_ram.memory\[511\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11564_ _04766_ _05171_ _05184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13972__B2 _05798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_168_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10786__A1 _04238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09640__A2 _03843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13303_ _06130_ _06401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_128_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10515_ _04469_ mod.u_cpu.rf_ram.memory\[440\]\[0\] _04470_ _04471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_11495_ _05128_ mod.u_cpu.rf_ram.memory\[284\]\[1\] _05136_ _05138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_14283_ _00137_ net3 mod.u_cpu.rf_ram.memory\[546\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_137_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07169__I _01477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13724__A1 _06382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09779__I0 _03936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13234_ _06280_ _06340_ _01197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10446_ _04422_ _00327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_196_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__15585__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_170_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10377_ _04363_ mod.u_cpu.rf_ram.memory\[462\]\[1\] _04374_ _04376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_13165_ _06273_ mod.u_cpu.rf_ram.memory\[349\]\[0\] _06274_ _06275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_156_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12116_ _05293_ _05471_ _05560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_13096_ _06217_ mod.u_cpu.rf_ram.memory\[59\]\[1\] _06231_ _06233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_151_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12047_ _05501_ mod.u_cpu.rf_ram.memory\[213\]\[1\] _05512_ _05514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_133_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_250_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_266_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_211_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_266_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07706__A2 mod.u_cpu.rf_ram.memory\[260\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08903__A1 _02527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_238_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13634__I _06455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_219_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_207_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13998_ mod.u_arbiter.i_wb_cpu_rdt\[12\] _06952_ _06958_ mod.u_arbiter.i_wb_cpu_dbus_dat\[12\]
+ _06961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_241_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_206_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12949_ mod.u_cpu.cpu.genblk1.align.ctrl_misal _06126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_248_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_209_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13570__S _06604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07565__S1 _01844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08762__S0 _02294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_179_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_261_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14619_ _00473_ net3 mod.u_cpu.rf_ram.memory\[378\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12186__S _05607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15599_ _01370_ net3 mod.u_cpu.rf_ram.memory\[120\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_53_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_221_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08140_ _01469_ _02281_ _02447_ _02448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__13963__A1 _03444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11813__I1 mod.u_cpu.rf_ram.memory\[49\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09092__B1 _03300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08071_ _02149_ _02364_ _02378_ _02379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__14802__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13015__I0 _06105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08985__A4 mod.u_cpu.cpu.state.o_cnt_r\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_31_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_259_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10529__A1 _04184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11577__I0 _05180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08198__A2 _02496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13191__A2 _03456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09294__I _03488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07945__A2 mod.u_cpu.rf_ram.memory\[238\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14952__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08973_ _03256_ _03277_ _03278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_69_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07924_ _01977_ _02187_ _02231_ _02232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_116_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_229_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07855_ _01819_ _02162_ _02163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_96_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15308__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_217_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_256_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_56_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07786_ mod.u_cpu.rf_ram.memory\[184\]\[0\] mod.u_cpu.rf_ram.memory\[185\]\[0\] mod.u_cpu.rf_ram.memory\[186\]\[0\]
+ mod.u_cpu.rf_ram.memory\[187\]\[0\] _02092_ _02093_ _02094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_227_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09525_ _03746_ _03747_ _03748_ _03749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_65_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_231_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_266_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__11501__I0 _05128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_225_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_213_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_225_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_197_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_213_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__14332__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_196_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09456_ _03365_ mod.u_cpu.cpu.bufreg.c_r _03680_ _03682_ _03683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__15458__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_197_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08407_ _02111_ _02713_ _02714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_36_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09387_ _03624_ _03620_ _03625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_184_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08338_ mod.u_cpu.rf_ram.memory\[509\]\[1\] _02645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_162_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09622__A2 _03829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14482__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07633__A1 _01938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08269_ _02551_ _02576_ _02577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_123_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_257_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10300_ _04298_ mod.u_cpu.rf_ram.memory\[474\]\[0\] _04323_ _04324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12509__A2 _05831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_193_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11280_ _04978_ mod.u_cpu.rf_ram.memory\[318\]\[0\] _04991_ _04992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_119_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13719__I _06320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10231_ _04274_ _00260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_180_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12623__I _05873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11193__A1 _04930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10162_ _03662_ _03753_ _04224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_126_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14970_ _00824_ net3 mod.u_cpu.rf_ram.memory\[57\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10093_ _04044_ _04174_ _04175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_121_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13921_ _06456_ _06468_ _06861_ _06452_ _06481_ _06899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_130_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_248_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_208_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13852_ _06842_ _06846_ _06483_ _06847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_75_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_223_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12803_ _06025_ _01081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_216_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13783_ _06739_ mod.u_arbiter.i_wb_cpu_rdt\[9\] _06455_ _06784_ _06785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_204_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10995_ _04794_ _00504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_188_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15522_ _01293_ net3 mod.u_cpu.cpu.immdec.imm19_12_20\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12734_ _05980_ _01057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_206_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_231_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09861__A2 _04014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_204_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14198__A1 _07076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_203_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15453_ _01227_ net3 mod.u_cpu.cpu.ctrl.o_ibus_adr\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__14825__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_203_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12665_ _05886_ _05934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_203_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_203_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12748__A2 _05422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14404_ _00258_ net3 mod.u_cpu.rf_ram.memory\[485\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11616_ _04539_ _05130_ _05218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_129_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15384_ _01159_ net3 mod.u_cpu.rf_ram.memory\[81\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_141_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12596_ _05888_ _05882_ _05889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_168_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14335_ _00189_ net3 mod.u_cpu.rf_ram.memory\[520\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11547_ _05159_ mod.u_cpu.rf_ram.memory\[275\]\[0\] _05172_ _05173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__11420__A2 _05085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_184_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_167_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14975__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_183_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14266_ _00120_ net3 mod.u_cpu.rf_ram.memory\[554\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_143_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11478_ _04852_ _05125_ _05126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_171_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13629__I _06332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13217_ _06321_ _06323_ _06324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13173__A2 _06140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10429_ _04411_ _00321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_152_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14197_ _07095_ _01405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_100_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07927__A2 _02234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12920__A2 _04704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13148_ mod.u_arbiter.i_wb_cpu_rdt\[25\] mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat\[9\]
+ _06263_ _06265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_152_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09047__C _03250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11149__I _04882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14122__A1 _03842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10053__I _03738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13079_ mod.u_cpu.rf_ram.memory\[105\]\[1\] _06221_ _06219_ _06222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09842__I _03994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08886__C _02465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12684__A1 _03895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_65_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11085__S _04856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_238_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07640_ _01643_ mod.u_cpu.rf_ram.memory\[292\]\[0\] _01947_ _01948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__14355__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07786__S1 _02093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07362__I _01669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_226_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15600__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_254_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07571_ _01710_ _01879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_213_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_207_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11813__S _05352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07538__S1 _01833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09310_ _03549_ _03559_ _03560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_178_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_22_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09241_ _03501_ _03502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13236__I0 _06273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_194_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09172_ mod.u_arbiter.i_wb_cpu_rdt\[14\] _03456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_187_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08123_ _02411_ _02430_ _02431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07615__A1 _01643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08126__C _02168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10228__I _03960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_257_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08054_ _02352_ _02355_ _02360_ _02361_ _02362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_190_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09368__A1 _03386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13164__A2 _04969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12443__I _03498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_227_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_157_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11175__A1 _04775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_115_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_248_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15130__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08591__A2 _02894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08956_ mod.u_arbiter.i_wb_cpu_dbus_we _03261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_4606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09752__I _03931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09915__I0 _04051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07907_ mod.u_cpu.rf_ram.memory\[209\]\[0\] _02215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_4639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3905 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08887_ _02455_ _03190_ _03193_ _02467_ _03194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_56_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13274__I _06371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3916 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10525__I1 mod.u_cpu.rf_ram.memory\[438\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3927 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_56_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3938 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07838_ _02104_ _02145_ _02146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_57_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3949 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15280__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_205_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_260_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12427__A1 _05019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14848__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07769_ _01677_ _02077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_112_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11723__S _05290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10289__I0 _04298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09508_ _03732_ _03733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_77_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10780_ _04569_ _04648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_52_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_72_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_198_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09439_ _03331_ _03670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_13_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_197_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__14998__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_185_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12450_ _05780_ mod.u_cpu.cpu.state.stage_two_req _05787_ _05788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_205_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_200_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11789__I0 _05329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11401_ _05069_ mod.u_cpu.rf_ram.memory\[2\]\[1\] _05072_ _05074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_122_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12381_ _05740_ _00944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_126_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14120_ _07041_ mod.u_cpu.rf_ram.memory\[11\]\[1\] _07044_ _07046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_166_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10461__I0 _04423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11332_ _05014_ mod.u_cpu.rf_ram.memory\[310\]\[1\] _05025_ _05027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_181_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07875__C _02164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14228__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_180_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_21_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09359__A1 _03489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14051_ _06914_ _07000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_84_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12353__I _05720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11263_ _04838_ _04969_ _04979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_137_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07909__A2 mod.u_cpu.rf_ram.memory\[208\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13002_ _06167_ _06164_ _06171_ _01134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_10214_ _03950_ _04262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08031__A1 _02090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11194_ _04918_ mod.u_cpu.rf_ram.memory\[331\]\[0\] _04931_ _04932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_121_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10913__A1 _01880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11961__I0 _05450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10145_ _04199_ mod.u_cpu.rf_ram.memory\[496\]\[1\] _04210_ _04212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_79_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_171_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14378__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_212_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15623__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_254_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_14953_ _00807_ net3 mod.u_cpu.rf_ram.memory\[529\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10076_ _04147_ _04162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12666__A1 _05896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13863__B1 _06837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09531__A1 _03754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08334__A2 mod.u_cpu.rf_ram.memory\[502\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13904_ _06707_ _06886_ _01321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10601__I _03713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08278__I _01636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14884_ _00738_ net3 mod.u_cpu.rf_ram.memory\[241\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_208_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07182__I mod.u_cpu.raddr\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_236_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_13835_ mod.u_cpu.cpu.immdec.imm7 _03682_ _06812_ _06831_ _06832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_169_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_250_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_216_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_13766_ mod.u_cpu.cpu.immdec.imm7 _06753_ _06769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_90_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_204_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10978_ mod.u_cpu.rf_ram.memory\[365\]\[1\] _04661_ _04781_ _04783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_71_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07910__I _01746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15505_ _01276_ net3 mod.u_arbiter.i_wb_cpu_dbus_adr\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_188_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12717_ _05969_ _01051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_189_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10249__S _04286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_189_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13697_ _06694_ _06431_ _06450_ _06705_ _06706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__15003__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13918__A1 _06451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_15436_ _01211_ net3 mod.u_cpu.rf_ram.memory\[91\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_129_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12648_ _05923_ mod.u_cpu.rf_ram.memory\[147\]\[1\] _05921_ _05924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_175_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_191_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15367_ _01142_ net3 mod.u_cpu.rf_ram.memory\[84\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12579_ _05877_ _01005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_102_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_200_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14318_ _00172_ net3 mod.u_cpu.rf_ram.memory\[528\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_171_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_15298_ _00058_ net4 mod.u_scanchain_local.module_data_in\[55\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_102_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15153__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12263__I _05634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14249_ _00103_ net3 mod.u_cpu.rf_ram.memory\[563\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_171_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11157__A1 _04360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07357__I _01499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08573__A2 _02879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08810_ mod.u_cpu.rf_ram.memory\[4\]\[1\] mod.u_cpu.rf_ram.memory\[5\]\[1\] mod.u_cpu.rf_ram.memory\[6\]\[1\]
+ mod.u_cpu.rf_ram.memory\[7\]\[1\] _02366_ _02383_ _03117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09790_ _03948_ _03961_ _03962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08741_ _01978_ _03038_ _03047_ _03048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09522__A1 _01850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08672_ mod.u_cpu.rf_ram.memory\[213\]\[1\] _02979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_187_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_253_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_242_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_214_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07623_ _01915_ _01917_ _01930_ _01812_ _01931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_54_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08089__A1 _02302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07554_ _01509_ _01862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13082__A1 _03932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09286__B1 _03536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_228_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07836__A1 _02124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07485_ mod.u_cpu.rf_ram.memory\[437\]\[0\] _01793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_195_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08137__B _02444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13909__A1 _06311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10691__I0 _04584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09224_ _03384_ _03486_ _03487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_158_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09155_ _03445_ _00009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_120_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_33_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09747__I _03733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08106_ _02410_ mod.u_cpu.rf_ram.memory\[22\]\[0\] _02413_ _01830_ _02414_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_163_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10443__I0 _04400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_162_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09086_ _03386_ _03387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_174_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08037_ _01493_ _02344_ _01534_ _02345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_107_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14520__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15646__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_190_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11943__I0 _05426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_249_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_231_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09988_ _04101_ _00190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_265_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_5148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_118_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_5159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_190_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_153_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_236_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08939_ _01464_ _01465_ _03206_ _03245_ _03246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XTAP_4425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14670__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08316__A2 mod.u_cpu.rf_ram.memory\[468\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11950_ _05450_ mod.u_cpu.rf_ram.memory\[21\]\[1\] _05447_ _05451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08098__I _01644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10123__A2 _03961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_218_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10901_ _04730_ _00474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_229_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11881_ _05262_ _05401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_232_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__15026__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13620_ _05164_ _04989_ _06636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10832_ _04682_ mod.u_cpu.rf_ram.memory\[388\]\[1\] _04680_ _04683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_72_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_198_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_198_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13551_ _06583_ _06594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_201_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10763_ _04626_ mod.u_cpu.rf_ram.memory\[3\]\[1\] _04634_ _04636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_158_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12671__I1 mod.u_cpu.rf_ram.memory\[121\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_186_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12502_ _05812_ _05827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_199_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10682__I0 _04579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13482_ _03602_ _06545_ _06546_ _03605_ _06548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_10694_ _04590_ _00407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_139_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15176__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15221_ _01074_ net3 mod.u_cpu.rf_ram.memory\[132\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12433_ _05642_ _05774_ _05775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07886__B _02193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11387__A1 _01964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_240_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15152_ _01005_ net3 mod.u_cpu.rf_ram.memory\[158\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_148_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12364_ _05710_ _05729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_181_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_14103_ _07028_ mod.u_cpu.rf_ram.memory\[110\]\[1\] _07033_ _07035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_11315_ _05015_ _00603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_15083_ _00937_ net3 mod.u_cpu.rf_ram.memory\[122\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12295_ _05677_ mod.u_cpu.rf_ram.memory\[188\]\[1\] _05680_ _05682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07177__I _01484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14034_ mod.u_arbiter.i_wb_cpu_rdt\[21\] _06987_ _06982_ mod.u_arbiter.i_wb_cpu_dbus_dat\[21\]
+ _06988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_11246_ _04967_ _00582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_49_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12887__A1 _05896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11934__I0 mod.u_cpu.rf_ram.memory\[169\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11177_ _04920_ _00560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_68_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10128_ _04200_ _00231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_255_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08307__A2 mod.u_cpu.rf_ram.memory\[476\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_209_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10331__I _04176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14936_ _00790_ net3 mod.u_cpu.rf_ram.memory\[224\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10059_ _04151_ _00211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_94_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_236_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07366__I0 mod.u_cpu.rf_ram.memory\[388\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4970 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_235_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4981 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_224_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4992 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_169_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14867_ _00721_ net3 mod.u_cpu.rf_ram.memory\[256\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_169_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_251_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11363__S _05048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13818_ _06814_ _06816_ _06817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_35_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13064__A1 _03918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14798_ _00652_ net3 mod.u_cpu.rf_ram.memory\[288\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_16_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12111__I0 _05539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_204_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08166__S1 _02473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13749_ _06335_ _03428_ _06754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_17_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15519__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_177_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07270_ _01560_ _01578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_149_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10673__I0 _04557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08491__A1 _01848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_192_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15419_ _01194_ net3 mod.u_cpu.rf_ram.memory\[349\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_258_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10425__I0 _04400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14543__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_89_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10506__I _04442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09991__A1 _03951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12178__I0 _05575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09911_ _04049_ _00165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_67_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_259_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14693__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_217_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08546__A2 _02844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09842_ _03994_ _04002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_98_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_247_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_218_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09773_ _03856_ _03939_ _03949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_67_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3009 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15049__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08724_ mod.u_cpu.rf_ram.memory\[245\]\[1\] _03031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__10241__I _03974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12350__I0 _05711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08655_ _02124_ _02954_ _02961_ _02143_ _02962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_214_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11853__A2 _03951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07606_ _01850_ _01914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08586_ _01978_ _02883_ _02892_ _02893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_241_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_230_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12102__I0 _05550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07550__I _01758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15199__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07537_ mod.u_cpu.rf_ram.memory\[336\]\[0\] mod.u_cpu.rf_ram.memory\[337\]\[0\] mod.u_cpu.rf_ram.memory\[338\]\[0\]
+ mod.u_cpu.rf_ram.memory\[339\]\[0\] _01843_ _01844_ _01845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_179_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11605__A2 _05210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_210_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07468_ _01774_ _01775_ _01776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_210_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_194_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09207_ _03476_ _00032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13358__A2 _06380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_183_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07399_ _01567_ _01706_ _01707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_124_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10416__I0 _04387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08381__I _01879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09138_ _03431_ _03387_ _03432_ _00074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_120_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10041__A1 _04044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09069_ _01433_ _03372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_190_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11100_ _03795_ _04868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_150_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12080_ _05535_ _05471_ _05536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_150_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_235_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11916__I0 _05426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10719__I1 mod.u_cpu.rf_ram.memory\[406\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11031_ mod.u_cpu.rf_ram.memory\[357\]\[1\] _04819_ _04816_ _04820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_81_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_237_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_264_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_218_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12097__A2 _05543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13294__A1 _06281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12982_ _06146_ _06155_ _06156_ _01129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_4266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_217_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_206_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14721_ _00575_ net3 mod.u_cpu.rf_ram.memory\[327\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_218_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11933_ _05078_ _05438_ _05439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_3554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14416__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_206_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14652_ _00506_ net3 mod.u_cpu.rf_ram.memory\[361\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11864_ _05385_ mod.u_cpu.rf_ram.memory\[70\]\[0\] _05389_ _05390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_17_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_127_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07460__I _01586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_233_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_13603_ mod.u_cpu.rf_ram.memory\[329\]\[1\] _06221_ _06621_ _06623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_2886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_242_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2897 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10815_ _04666_ mod.u_cpu.rf_ram.memory\[391\]\[1\] _04670_ _04672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__13597__A2 _03694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_14_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14583_ _00437_ net3 mod.u_cpu.rf_ram.memory\[396\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11795_ _05341_ _00757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_159_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_198_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10655__I0 _04560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14566__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13534_ mod.u_arbiter.i_wb_cpu_dbus_adr\[2\] mod.u_arbiter.i_wb_cpu_dbus_adr\[3\]
+ _06584_ _06585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_207_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_201_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10746_ _04625_ _00424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_41_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10280__A1 _04307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_186_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13349__A2 _06445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13465_ _06536_ _01232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_145_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10677_ _04579_ mod.u_cpu.rf_ram.memory\[414\]\[1\] _04576_ _04580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_199_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15204_ _01057_ net3 mod.u_cpu.rf_ram.memory\[136\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_145_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12416_ mod.u_cpu.rf_ram.memory\[489\]\[0\] _05622_ _05763_ _05764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_13396_ _06483_ _06489_ _06490_ _06491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_126_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08776__A2 _03082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11080__I0 _04841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15135_ _00988_ net3 mod.u_cpu.rf_ram.memory\[469\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_142_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12347_ _04014_ _05703_ _05717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_86_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15066_ _00920_ net3 mod.u_cpu.rf_ram.memory\[186\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12278_ _05660_ mod.u_cpu.rf_ram.memory\[191\]\[1\] _05669_ _05671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__11907__I0 _05406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14017_ mod.u_arbiter.i_wb_cpu_dbus_dat\[18\] _06966_ _06975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11229_ _04107_ _04955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__08084__S0 _02391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_214_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12580__I0 _05874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13285__A1 _06367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_95_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_224_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10996__I _03761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12189__S _05607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14919_ _00773_ net3 mod.u_cpu.rf_ram.memory\[159\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__15341__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13372__I _06292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08700__A2 mod.u_cpu.rf_ram.memory\[198\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08440_ _02143_ _02744_ _02746_ _02747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__10894__I0 _04695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_224_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_223_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__14909__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_212_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07370__I _01677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08839__I0 _03142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08371_ _02665_ _02667_ _02676_ _02677_ _02678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_56_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_225_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_177_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07322_ _01490_ _01630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08464__A1 _02059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15491__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07267__A2 _01574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_176_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_220_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07253_ _01560_ _01561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_176_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12399__I0 _05745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_192_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07184_ _01491_ _01492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_129_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08134__C _02166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_191_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_254_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07973__C _02280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_232_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_160_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_235_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12571__I0 _05869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09825_ _03988_ _00140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_63_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14439__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_219_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__11067__I _04844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_246_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09756_ _03935_ _00124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_58_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12323__I0 _05696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08707_ _02385_ mod.u_cpu.rf_ram.memory\[236\]\[1\] _03014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_55_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09687_ _03877_ mod.u_cpu.rf_ram.memory\[55\]\[0\] _03880_ _03881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__11826__A2 _03942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_104_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_266_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_265_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14589__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08638_ mod.u_cpu.rf_ram.memory\[168\]\[1\] mod.u_cpu.rf_ram.memory\[169\]\[1\] mod.u_cpu.rf_ram.memory\[170\]\[1\]
+ mod.u_cpu.rf_ram.memory\[171\]\[1\] _02106_ _02127_ _02945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_203_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_199_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08569_ mod.u_cpu.rf_ram.memory\[277\]\[1\] _02876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_70_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10600_ _04526_ _00377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07258__A2 _01555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08455__A1 _01496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11580_ _05194_ mod.u_cpu.rf_ram.memory\[270\]\[1\] _05192_ _05195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_161_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09201__S _03469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_211_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10531_ _01793_ _04479_ _04480_ _00354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_195_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13250_ _06350_ _01203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13200__A1 _06283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10462_ _04433_ _00332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_108_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12201_ mod.u_cpu.rf_ram.memory\[201\]\[1\] _05617_ _05615_ _05618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_129_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_202_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__13751__A2 _06425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_13181_ _06286_ _06287_ _06288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_129_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10393_ _04387_ mod.u_cpu.rf_ram.memory\[460\]\[1\] _04385_ _04388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_109_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_191_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10565__A2 _04447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15214__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12132_ _05566_ mod.u_cpu.rf_ram.memory\[208\]\[1\] _05569_ _05571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_135_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11178__S _04919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09707__A1 _03893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13457__I _06513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12063_ _04983_ _03771_ _05525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_172_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10082__S _04165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07455__I _01762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09871__S _04020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11014_ _04250_ _04808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_150_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15364__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4030 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_265_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4041 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4052 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_161_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4063 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4074 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4085 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_161_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12965_ _06135_ _06141_ _01127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_206_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4096 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11705__I _05262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11916_ _05426_ mod.u_cpu.rf_ram.memory\[223\]\[1\] _05424_ _05427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_14704_ _00558_ net3 mod.u_cpu.rf_ram.memory\[335\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_46_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08286__I _02116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07497__A2 mod.u_cpu.rf_ram.memory\[444\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_205_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12896_ _06086_ mod.u_cpu.rf_ram.memory\[98\]\[1\] _06084_ _06087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07190__I _01497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_260_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_221_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_221_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14635_ _00489_ net3 mod.u_cpu.rf_ram.memory\[370\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_178_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11847_ _05377_ _00773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07123__C _01431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1960 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1971 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10628__I0 _04537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1982 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14566_ _00420_ net3 mod.u_cpu.rf_ram.memory\[404\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1993 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08446__A1 _02730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11778_ _05330_ _00751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12242__A2 _05611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_201_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08836__I3 mod.u_cpu.rf_ram.memory\[51\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13517_ _03425_ _06570_ _06571_ _01249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_202_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10729_ _04613_ _00419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_119_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14497_ _00351_ net3 mod.u_cpu.rf_ram.memory\[43\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_105_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_220_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_13448_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[8\] _06525_ _06526_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[9\]
+ _06527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__13042__I1 mod.u_cpu.rf_ram.memory\[107\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10005__A1 _03961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09946__A1 _03886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13742__A2 _06712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13379_ _06454_ _06475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_154_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11753__A1 _05312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_170_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15118_ _00971_ net3 mod.u_cpu.rf_ram.memory\[449\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_255_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_255_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_114_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15049_ _00903_ net3 mod.u_cpu.rf_ram.memory\[195\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_07940_ _02244_ mod.u_cpu.rf_ram.memory\[236\]\[0\] _02247_ _02248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07972__A3 _02279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_218_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11505__A1 _04868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07365__I _01672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_229_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07871_ _01646_ _02179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10859__A3 _03724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_256_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09610_ _03746_ _03819_ _03820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_228_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08921__A2 _03227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13258__A1 _03390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14731__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09580__I _03795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09541_ _03763_ _03764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_97_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_252_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09721__I1 mod.u_cpu.rf_ram.memory\[556\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09472_ _03697_ _03698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_64_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_262_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_08423_ _01914_ _02730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_224_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_251_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14881__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_240_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08354_ _02654_ _02655_ _02659_ _02660_ _02661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__08437__A1 _01680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07968__C _01766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_220_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07305_ _01578_ _01612_ _01613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12446__I _05783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08988__A2 _03292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08285_ _02591_ _02592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_177_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11992__A1 _03767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15237__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07236_ _01508_ mod.u_cpu.rf_ram.memory\[460\]\[0\] _01543_ _01544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_153_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13033__I1 mod.u_cpu.rf_ram.memory\[108\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07167_ _01469_ _01471_ _01475_ _01476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_173_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11744__A1 _04983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_191_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14261__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15387__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_259_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12544__I0 _05837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09808_ _03948_ _03975_ _03976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_189_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_247_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_228_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09739_ _03890_ mod.u_cpu.rf_ram.memory\[554\]\[1\] _03920_ _03922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_216_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12750_ _02162_ _05989_ _05990_ _01063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__09712__I1 _03735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08676__A1 _01705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_242_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_188_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_216_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11701_ _05268_ mod.u_cpu.rf_ram.memory\[252\]\[0\] _05276_ _05277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_37_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10483__A1 _04439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_152_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08771__S1 _02323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12681_ _05945_ _01039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14420_ _00274_ net3 mod.u_cpu.rf_ram.memory\[477\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_230_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11632_ _03733_ _05229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08428__A1 _02526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12224__A2 _05632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07878__C _02185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14351_ _00205_ net3 mod.u_cpu.rf_ram.memory\[512\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11563_ _05183_ _00683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_211_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_168_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13302_ _06366_ _06376_ _06381_ _06399_ _06400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_156_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10514_ _04168_ _04464_ _04470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_14282_ _00136_ net3 mod.u_cpu.rf_ram.memory\[546\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11494_ _05137_ _00660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_196_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14604__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13233_ _06325_ _06333_ _06336_ _06339_ _06340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_137_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13724__A2 _06493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10445_ _04410_ mod.u_cpu.rf_ram.memory\[451\]\[1\] _04420_ _04422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_109_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08600__A1 _02136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13164_ _05515_ _04969_ _06274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10376_ _04375_ _00304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_151_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_237_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__13187__I _06284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12091__I _05387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12115_ _05520_ _05559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_13095_ _06232_ _01166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_112_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07185__I _01492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14754__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12046_ _02226_ _05512_ _05513_ _00836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_49_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_215_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_238_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__12160__A1 _05588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_65_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_266_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_226_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13997_ mod.u_arbiter.i_wb_cpu_dbus_dat\[13\] _06954_ _06960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_207_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07134__B _01441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_234_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_207_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12948_ _06122_ _06123_ _06124_ _06125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_3170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_207_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_261_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_222_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08762__S1 _02295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_233_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12879_ _06070_ mod.u_cpu.rf_ram.memory\[246\]\[1\] _06074_ _06076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_2480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08419__A1 _02534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14618_ _00472_ net3 mod.u_cpu.rf_ram.memory\[378\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__13412__A1 _03910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15598_ _01369_ net3 mod.u_cpu.rf_ram.memory\[120\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_261_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_187_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11274__I0 _04976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14549_ _00403_ net3 mod.u_cpu.rf_ram.memory\[413\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12266__I _05604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_222_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_202_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09092__A1 _03362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_179_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09092__B2 _03279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11974__A1 _03893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08070_ _02365_ _02368_ _02376_ _02377_ _02378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_174_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14284__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11726__A1 _05293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10529__A2 _04447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11577__I1 mod.u_cpu.rf_ram.memory\[270\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12774__I0 mod.u_cpu.rf_ram.memory\[133\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08412__C _01992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08972_ _03268_ _03270_ _03276_ _03277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_130_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07923_ _02195_ _02208_ _02229_ _02230_ _01978_ _02231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_190_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_257_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07854_ mod.u_cpu.rf_ram.memory\[199\]\[0\] _02162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_28_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_229_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10701__A2 _03933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07785_ _02042_ _02093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09524_ _03709_ _03748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_266_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08658__A1 _02944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_213_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13651__A1 _06661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_224_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_149_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10465__A1 _03755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09455_ _03349_ _03681_ _03682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_101_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_51_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13560__I _06583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_213_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_213_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_197_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08406_ mod.u_cpu.rf_ram.memory\[445\]\[1\] _02713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_212_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13403__A1 _06432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09386_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[25\] _03624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07698__C _02005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_178_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_212_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__14627__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_196_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08337_ mod.u_cpu.rf_ram.memory\[504\]\[1\] mod.u_cpu.rf_ram.memory\[505\]\[1\] mod.u_cpu.rf_ram.memory\[506\]\[1\]
+ mod.u_cpu.rf_ram.memory\[507\]\[1\] _02385_ _02633_ _02644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_123_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_193_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07633__A2 mod.u_cpu.rf_ram.memory\[310\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08830__A1 _02410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08268_ mod.u_cpu.rf_ram.memory\[543\]\[0\] _02576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_126_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_193_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_203_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_193_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07219_ _01490_ _01527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_152_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12904__I _05720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08199_ _02209_ _02507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_152_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_192_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_152_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08603__B _02046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14777__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10230_ _04249_ mod.u_cpu.rf_ram.memory\[484\]\[0\] _04273_ _04274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_69_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_238_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10161_ _04222_ _04223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_134_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09138__A2 _03387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10092_ _04172_ _04173_ _04174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_266_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13920_ _06898_ _01325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_120_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08897__A1 _02471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07733__I _01743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13851_ _06451_ _06672_ _06844_ _06845_ _06846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_142_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11255__I _04125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_12802_ _06010_ mod.u_cpu.rf_ram.memory\[128\]\[0\] _06024_ _06025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_13782_ _03509_ mod.u_arbiter.i_wb_cpu_rdt\[25\] _06784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__15402__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10994_ _04774_ mod.u_cpu.rf_ram.memory\[362\]\[0\] _04793_ _04794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_43_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_262_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_243_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15521_ _01292_ net3 mod.u_cpu.cpu.immdec.imm19_12_20\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12733_ _05963_ mod.u_cpu.rf_ram.memory\[136\]\[0\] _05979_ _05980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_204_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_215_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_204_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07321__A1 _01602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_16_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15452_ _01226_ net3 mod.u_cpu.cpu.ctrl.o_ibus_adr\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_76_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12664_ _05933_ _01034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_188_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_231_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_243_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14403_ _00257_ net3 mod.u_cpu.rf_ram.memory\[486\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11615_ _05217_ _00701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_89_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_204_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15552__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15383_ _01158_ net3 mod.u_cpu.rf_ram.memory\[81\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_184_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12595_ _03789_ _05888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_196_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14334_ _00188_ net3 mod.u_cpu.rf_ram.memory\[520\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11546_ _05037_ _05171_ _05172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_156_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_204_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08821__A1 _02410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14265_ _00119_ net3 mod.u_cpu.rf_ram.memory\[555\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11477_ _05124_ _05125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_137_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13216_ _06322_ _06323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_48_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10428_ _04410_ mod.u_cpu.rf_ram.memory\[454\]\[1\] _04408_ _04411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_174_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14196_ _06057_ _03388_ _07095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_124_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08232__C _02539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13147_ _06264_ _01186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10359_ _04363_ mod.u_cpu.rf_ram.memory\[465\]\[1\] _04361_ _04364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14122__A2 _05631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13078_ _03734_ _06221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_250_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_266_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_239_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11366__S _05048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12029_ _05239_ _03851_ _05503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_22_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08888__A1 _02449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12684__A2 _05589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13881__A1 _06426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_266_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10695__A1 _04322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07560__A1 _01863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07570_ _01875_ mod.u_cpu.rf_ram.memory\[372\]\[0\] _01877_ _01878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_53_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15082__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_206_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_146_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_234_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_222_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11495__I0 _05128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07312__A1 _01592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_181_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09240_ _03500_ _03501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_61_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_210_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_210_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11247__I0 _04952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13397__B1 _06481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_221_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_178_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09171_ _03455_ _00015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07311__C _01618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09065__A1 _03300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08112__I0 mod.u_cpu.rf_ram.memory\[52\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11947__A1 _05448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08122_ mod.u_cpu.rf_ram.memory\[39\]\[0\] _02430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_147_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_222_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07615__A2 mod.u_cpu.rf_ram.memory\[316\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08053_ _01528_ _02361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07818__I _01568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11175__A2 _04906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_5308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08955_ mod.u_cpu.cpu.state.o_cnt_r\[0\] _03259_ _03260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07981__C _02139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_233_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07906_ _02209_ _02210_ _02213_ _02214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_57_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_243_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08886_ _02461_ mod.u_cpu.rf_ram.memory\[574\]\[1\] _03192_ _02465_ _03193_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_29_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13872__A1 _03503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15425__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3906 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_217_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3917 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_256_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3928 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07837_ _02105_ _02123_ _02144_ _02145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_110_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3939 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_186_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12427__A2 _04442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07768_ _02074_ _02075_ _01602_ _02076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_244_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_225_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09507_ _01462_ _03352_ _03731_ _03732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_225_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__10289__I1 mod.u_cpu.rf_ram.memory\[476\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15575__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07699_ _01787_ _02007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__07303__A1 _01607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_213_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09438_ _03668_ _03669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_12_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_160_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_185_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_184_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09369_ _03568_ _03607_ _03608_ _03609_ _00064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_197_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_240_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_201_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11400_ _05073_ _00630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08803__A1 _02190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12380_ _05731_ mod.u_cpu.rf_ram.memory\[178\]\[0\] _05739_ _05740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_123_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11331_ _05026_ _00608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_115_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_158_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14050_ _06997_ _06999_ _01354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_125_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11262_ _04960_ _04978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_180_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08052__C _02359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13001_ mod.u_cpu.cpu.genblk3.csr.mcause3_0\[3\] _03353_ _06163_ _06170_ _06171_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_238_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10213_ _04261_ _00255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10154__I _03885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11193_ _04930_ _04926_ _04931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_106_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10144_ _04211_ _00236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_251_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14952_ _00806_ net3 mod.u_cpu.rf_ram.memory\[529\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_130_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10075_ _04161_ _00217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_248_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12666__A2 _05721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13863__B2 mod.u_cpu.cpu.immdec.imm24_20\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07463__I _01569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09531__A2 _03721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13903_ _03355_ _06140_ _06886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_14883_ _00737_ net3 mod.u_cpu.rf_ram.memory\[242\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_35_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_210_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_13834_ _06651_ _06829_ _06830_ _03682_ _06831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__13615__A1 _04844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_249_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_204_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13765_ _06768_ _01300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10977_ _01894_ _04781_ _04782_ _00498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_15_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_188_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15504_ _01275_ net3 mod.u_arbiter.i_wb_cpu_dbus_adr\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12716_ _05963_ mod.u_cpu.rf_ram.memory\[138\]\[0\] _05968_ _05969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__14942__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13696_ _06295_ _06306_ _06464_ _06682_ _06493_ _06323_ _06705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_203_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_15435_ _01210_ net3 mod.u_cpu.cpu.immdec.imm11_7\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12647_ _05873_ _05923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09047__A1 _03349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14040__A1 mod.u_arbiter.i_wb_cpu_dbus_dat\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_200_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15366_ _01141_ net3 mod.u_cpu.rf_ram.memory\[10\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_156_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_200_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12578_ _05869_ mod.u_cpu.rf_ram.memory\[158\]\[0\] _05876_ _05877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_172_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_190_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11529_ _05159_ mod.u_cpu.rf_ram.memory\[278\]\[0\] _05160_ _05161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_14317_ _00171_ net3 mod.u_cpu.rf_ram.memory\[52\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_129_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15297_ _00057_ net4 mod.u_scanchain_local.module_data_in\[54\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12729__I0 _05966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14248_ _00102_ net3 mod.u_cpu.rf_ram.memory\[563\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_132_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_217_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11157__A2 _04906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12354__A1 _05452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__13576__S _06604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11401__I0 _05069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14179_ _07084_ _01398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__14322__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_140_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15448__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08897__C _02518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11096__S _04865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13375__I _06470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12106__A1 _05488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07781__A1 _01818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08740_ _03017_ _03039_ _03046_ _01870_ _03047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_39_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13854__A1 _06847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08405__S0 _02711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07373__I _01509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_238_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_227_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08671_ _02606_ _02977_ _02978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__14472__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_266_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_227_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15598__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11824__S _05359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07622_ _01918_ _01923_ _01928_ _01929_ _01930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_93_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_254_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_199_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_226_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_207_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07553_ _01857_ mod.u_cpu.rf_ram.memory\[380\]\[0\] _01860_ _01861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08089__A2 mod.u_cpu.rf_ram.memory\[28\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09286__A1 _03535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13082__A2 _06223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07836__A2 _02128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07484_ mod.u_cpu.rf_ram.memory\[432\]\[0\] mod.u_cpu.rf_ram.memory\[433\]\[0\] mod.u_cpu.rf_ram.memory\[434\]\[0\]
+ mod.u_cpu.rf_ram.memory\[435\]\[0\] _01745_ _01747_ _01792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_107_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_263_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_250_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_210_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08137__C _01591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09223_ _03406_ _03486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_166_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10840__A1 _04281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_179_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_210_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09154_ mod.u_arbiter.i_wb_cpu_rdt\[7\] _03444_ _03442_ _03445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09589__A2 _03786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_175_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08105_ _02411_ _02412_ _02413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_148_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11640__I0 _05234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10443__I1 mod.u_cpu.rf_ram.memory\[451\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09085_ _03385_ _03386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08261__A2 mod.u_cpu.rf_ram.memory\[534\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07548__I _01603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08036_ mod.u_cpu.rf_ram.memory\[92\]\[0\] mod.u_cpu.rf_ram.memory\[93\]\[0\] mod.u_cpu.rf_ram.memory\[94\]\[0\]
+ mod.u_cpu.rf_ram.memory\[95\]\[0\] _01636_ _01638_ _02344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_123_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_192_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_192_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09987_ _04096_ mod.u_cpu.rf_ram.memory\[51\]\[0\] _04100_ _04101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_5127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14815__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08600__C _01504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_258_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08938_ _01459_ _03225_ _03244_ _03245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XTAP_4415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_218_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_257_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08869_ _02542_ _03168_ _03175_ _02518_ _03176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_3725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11734__S _05297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10900_ _04728_ mod.u_cpu.rf_ram.memory\[377\]\[0\] _04729_ _04730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_3758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_260_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11880_ _05400_ _00783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__14965__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_233_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09204__S _03474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10831_ _04640_ _04682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_72_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13550_ _06593_ _01260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_10762_ _04635_ _00430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_13_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09003__I mod.u_cpu.cpu.alu.i_rs1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12501_ _05826_ _00978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_185_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_232_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_186_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13481_ _06547_ _01237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_240_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_185_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10693_ _04579_ mod.u_cpu.rf_ram.memory\[411\]\[1\] _04588_ _04590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_157_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09938__I _04067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15220_ _01073_ net3 mod.u_cpu.rf_ram.memory\[132\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12432_ _05593_ _05438_ _05774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_201_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07886__C _01666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15151_ _01004_ net3 mod.u_cpu.rf_ram.memory\[15\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_154_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12363_ _05728_ _00938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_181_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__14345__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07458__I _01765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14102_ _07034_ _01371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_11314_ _05014_ mod.u_cpu.rf_ram.memory\[313\]\[1\] _05012_ _05015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_154_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_15082_ _00936_ net3 mod.u_cpu.rf_ram.memory\[122\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12294_ _05681_ _00916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_154_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14033_ _06963_ _06987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_101_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11245_ _04961_ mod.u_cpu.rf_ram.memory\[323\]\[0\] _04966_ _04967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_106_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_141_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12887__A2 _06080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11934__I1 _05437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11176_ _04918_ mod.u_cpu.rf_ram.memory\[334\]\[0\] _04919_ _04920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_45_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14495__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10127_ _04199_ mod.u_cpu.rf_ram.memory\[4\]\[1\] _04197_ _04200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_110_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_249_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_236_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_94_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14935_ _00789_ net3 mod.u_cpu.rf_ram.memory\[225\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11698__I0 _05271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10058_ _04140_ mod.u_cpu.rf_ram.memory\[50\]\[1\] _04149_ _04151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_209_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4960 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4971 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_169_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_247_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4982 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_180_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_236_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_180_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4993 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14866_ _00720_ net3 mod.u_cpu.rf_ram.memory\[256\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_208_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_250_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_236_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_169_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13817_ _06423_ _06449_ _06459_ _06816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_63_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14797_ _00651_ net3 mod.u_cpu.rf_ram.memory\[28\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_51_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13064__A2 _06092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12111__I1 mod.u_cpu.rf_ram.memory\[68\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_189_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13748_ _06482_ _06753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_148_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10673__I1 mod.u_cpu.rf_ram.memory\[414\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__15120__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13679_ mod.u_cpu.cpu.immdec.imm19_12_20\[2\] _06678_ _06690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08491__A2 _02777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15418_ _01193_ net3 mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_78_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_191_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10425__I1 mod.u_cpu.rf_ram.memory\[454\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12274__I _05667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15349_ _01124_ net3 mod.u_cpu.rf_ram.memory\[369\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__15270__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14838__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12178__I1 mod.u_cpu.rf_ram.memory\[204\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09910_ _04036_ mod.u_cpu.rf_ram.memory\[532\]\[1\] _04047_ _04049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_132_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10889__A1 _04414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09841_ _03915_ _04001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_28_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_224_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08199__I _02209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09772_ _03766_ _03948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_140_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14988__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08723_ mod.u_cpu.rf_ram.memory\[240\]\[1\] mod.u_cpu.rf_ram.memory\[241\]\[1\] mod.u_cpu.rf_ram.memory\[242\]\[1\]
+ mod.u_cpu.rf_ram.memory\[243\]\[1\] _01647_ _01732_ _03030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_100_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_239_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07506__A1 _01791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_227_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_227_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08654_ _02110_ _02957_ _02960_ _02141_ _02961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_2309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_242_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_255_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_199_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_187_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07831__I _01746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07605_ _01835_ _01847_ _01912_ _01482_ _01913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_26_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_199_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08585_ _01992_ _02884_ _02891_ _02007_ _02892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__12449__I _05786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07536_ _01503_ _01844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_81_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_223_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_167_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_222_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_167_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07467_ mod.u_cpu.rf_ram.memory\[429\]\[0\] _01775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_161_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14368__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09206_ mod.u_arbiter.i_wb_cpu_rdt\[28\] mod.u_arbiter.i_wb_cpu_dbus_dat\[25\] _03474_
+ _03476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_202_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15613__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07398_ mod.u_cpu.rf_ram.memory\[413\]\[0\] _01706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_124_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__12184__I _03909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13763__B1 _06765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10416__I1 mod.u_cpu.rf_ram.memory\[456\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09137_ mod.u_arbiter.i_wb_cpu_rdt\[3\] _03410_ _03432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_147_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_194_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09068_ mod.u_arbiter.i_wb_cpu_ibus_adr\[0\] _03371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_190_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07993__A1 _02297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11729__S _05294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08019_ _02298_ _02326_ _02327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_78_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10633__S _04548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_190_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08617__S0 _02022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08611__B _01662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11030_ _04531_ _04819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_249_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13118__I0 _06237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_265_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10432__I _03898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_77_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_134_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_182_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12981_ mod.u_cpu.cpu.genblk3.csr.mie_mtie _06155_ _06056_ _06156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_4256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_218_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13294__A2 _06284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14720_ _00574_ net3 mod.u_cpu.rf_ram.memory\[327\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_218_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11932_ _03892_ _05319_ _05438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__09442__B _03669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_261_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10352__I0 _04345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_232_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_233_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11863_ _05355_ _05388_ _05389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_166_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14651_ _00505_ net3 mod.u_cpu.rf_ram.memory\[362\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__15143__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12359__I _05666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_214_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13602_ _06622_ _01283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09869__S _04020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10814_ _04671_ _00446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2898 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10104__I0 _04178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11794_ mod.u_cpu.rf_ram.memory\[233\]\[1\] _05230_ _05339_ _05341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_220_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_198_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14582_ _00436_ net3 mod.u_cpu.rf_ram.memory\[396\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10804__A1 _04255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10745_ _04622_ mod.u_cpu.rf_ram.memory\[402\]\[0\] _04624_ _04625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_41_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13533_ _06583_ _06584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_185_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09668__I _03865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15293__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13464_ _03574_ _06531_ _06532_ _03578_ _06536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_10676_ _04578_ _04579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_186_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_173_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15203_ _01056_ net3 mod.u_cpu.rf_ram.memory\[78\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_145_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12415_ _05588_ _04228_ _05763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__10607__I _04531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13395_ _06310_ _06329_ _06490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_126_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08076__I2 mod.u_cpu.rf_ram.memory\[6\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_12346_ _05716_ _00933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_15134_ _00987_ net3 mod.u_cpu.rf_ram.memory\[469\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_177_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07984__A1 _02124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15065_ _00919_ net3 mod.u_cpu.rf_ram.memory\[187\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12822__I _06018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12277_ _05670_ _00910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_114_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08608__S0 _02638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14016_ _06973_ _06974_ _01345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_218_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11228_ _03924_ _04954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_136_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08084__S1 _01720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_229_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10342__I _03850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11159_ _04908_ _00554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_96_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13809__A1 _06401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_191_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_255_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_209_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13285__A2 _06382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09352__B _03488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14918_ _00772_ net3 mod.u_cpu.rf_ram.memory\[159\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_237_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_224_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_4790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_184_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_75_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_251_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14849_ _00703_ net3 mod.u_cpu.rf_ram.memory\[263\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_91_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_224_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11048__A1 _04831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08370_ _01886_ _02677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_56_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14510__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15636__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08839__I1 _03143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_205_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12796__A1 _05870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07321_ _01602_ _01621_ _01628_ _01587_ _01629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_204_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_149_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_221_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08464__A2 mod.u_cpu.rf_ram.memory\[372\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07252_ mod.u_cpu.raddr\[0\] _01560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_143_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14660__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07183_ _01490_ _01491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08847__S0 _01647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_219_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_160_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15016__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07826__I _01634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12020__I0 _05484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_193_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_98_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07727__A1 _01977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11348__I _04989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_247_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12571__I1 mod.u_cpu.rf_ram.memory\[15\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09824_ _03958_ mod.u_cpu.rf_ram.memory\[544\]\[0\] _03987_ _03988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_86_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10582__I0 _04514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_228_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09755_ _03916_ mod.u_cpu.rf_ram.memory\[552\]\[0\] _03934_ _03935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_39_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15166__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09024__S0 mod.u_cpu.cpu.bufreg.lsb\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12323__I1 mod.u_cpu.rf_ram.memory\[179\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11287__A1 _04994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08706_ mod.u_cpu.rf_ram.memory\[237\]\[1\] _03013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_73_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_251_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_230_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09686_ _03878_ _03879_ _03880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_243_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_214_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08152__A1 _02456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_215_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08637_ _02938_ _02943_ _02102_ _02944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_215_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_230_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12087__I0 _05539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09689__S _03880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08568_ mod.u_cpu.rf_ram.memory\[272\]\[1\] mod.u_cpu.rf_ram.memory\[273\]\[1\] mod.u_cpu.rf_ram.memory\[274\]\[1\]
+ mod.u_cpu.rf_ram.memory\[275\]\[1\] _01957_ _01958_ _02875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_202_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07519_ _01700_ _01827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_120_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08499_ _02668_ _02802_ _02805_ _02096_ _02806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_22_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08455__A2 mod.u_cpu.rf_ram.memory\[380\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_195_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09488__I _03713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_195_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10530_ _04439_ _04479_ _04480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_196_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10262__A2 _04295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_183_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13736__B1 _06741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10461_ _04423_ mod.u_cpu.rf_ram.memory\[448\]\[0\] _04432_ _04433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_183_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09404__A1 mod.u_arbiter.i_wb_cpu_dbus_adr\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08838__S0 _02242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13200__A2 _06285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_182_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12200_ _05229_ _05617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_136_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13180_ _05783_ mod.u_arbiter.i_wb_cpu_rdt\[12\] _06287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_135_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10392_ _04344_ _04387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_109_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_164_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07966__A1 _02180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12131_ _05570_ _00864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_151_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12642__I _05372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_12062_ _05524_ _00841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09707__A2 _03896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15509__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11013_ _04807_ _00509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_89_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10573__I0 _04506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_237_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08391__A1 _02191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15821_ net4 net6 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_4020 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_219_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4031 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4042 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4053 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_4064 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_161_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_248_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_219_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_206_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4075 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_161_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_219_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4086 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12964_ mod.u_cpu.cpu.ctrl.i_iscomp _06140_ _06141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__14533__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_218_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07471__I _01778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4097 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_233_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14703_ _00557_ net3 mod.u_cpu.rf_ram.memory\[336\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_79_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11915_ _05405_ _05426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_206_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12895_ _06018_ _06086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_2651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_206_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14634_ _00488_ net3 mod.u_cpu.rf_ram.memory\[370\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_57_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11846_ _05364_ mod.u_cpu.rf_ram.memory\[159\]\[1\] _05375_ _05377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_2684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_221_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1950 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_221_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_207_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1961 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1972 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14683__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1983 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10628__I1 mod.u_cpu.rf_ram.memory\[422\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13422__B net5 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11777_ _05329_ mod.u_cpu.rf_ram.memory\[236\]\[1\] _05326_ _05330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_202_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14565_ _00419_ net3 mod.u_cpu.rf_ram.memory\[405\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08446__A2 _02752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_207_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1994 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10728_ _04608_ mod.u_cpu.rf_ram.memory\[405\]\[1\] _04610_ _04613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_13516_ _03426_ _06570_ _06571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_186_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14496_ _00350_ net3 mod.u_cpu.rf_ram.memory\[43\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_173_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10659_ _04566_ _00396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_13447_ _06513_ _06526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__15039__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13378_ _06462_ _06467_ _06469_ _06473_ _06474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_115_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12950__A1 _06116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_182_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15117_ _00970_ net3 mod.u_cpu.rf_ram.memory\[519\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_177_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12329_ _05696_ mod.u_cpu.rf_ram.memory\[184\]\[0\] _05704_ _05705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_142_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12002__I0 _05484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15048_ _00902_ net3 mod.u_cpu.rf_ram.memory\[195\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_141_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15189__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07709__A1 _01722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12702__A1 _03728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_190_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07870_ _02175_ mod.u_cpu.rf_ram.memory\[204\]\[0\] _02177_ _02178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_69_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_205_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13258__A2 _03672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09540_ _03762_ _03763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_110_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_237_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10800__I _04531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08134__A1 _02155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07381__I _01633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtiny_user_project_180 wbs_dat_o[30] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_92_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09471_ _03696_ _03697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_225_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__14207__A1 _03895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_1243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09882__A1 _03805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_212_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08422_ _02692_ mod.u_cpu.rf_ram.memory\[414\]\[1\] _02728_ _01773_ _02729_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_110_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12069__I0 _05521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_225_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_211_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13332__B _06330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08353_ _01679_ _02660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_177_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08437__A2 _02743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08288__I2 mod.u_cpu.rf_ram.memory\[458\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07304_ mod.u_cpu.rf_ram.memory\[511\]\[0\] _01612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_71_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08284_ _01851_ _02591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09101__I _03401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_260_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11992__A2 _04026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07235_ _01511_ _01542_ _01543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_192_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10247__I _04125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07166_ _01474_ _01475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_180_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07984__C _02291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14406__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07948__A1 _01740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11744__A2 _03823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07556__I _01671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_191_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_232_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14556__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_219_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08373__A1 _01591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_189_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09807_ _03974_ _03975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__13507__B _06562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07999_ _02302_ mod.u_cpu.rf_ram.memory\[110\]\[0\] _02305_ _02306_ _02307_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_87_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_262_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09738_ _03921_ _00120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_132_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__10307__I0 _04326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_216_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08125__A1 _02405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_215_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09173__I0 _03456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_216_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09669_ _03855_ _03866_ _03867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08676__A2 _02982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11742__S _05302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_231_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11700_ _04859_ _05255_ _05276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_199_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_167_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12680_ _05934_ mod.u_cpu.rf_ram.memory\[142\]\[0\] _05944_ _05945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_1246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_203_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11631_ _02012_ _05227_ _05228_ _00706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_145_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08428__A2 _02734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11562_ _05178_ mod.u_cpu.rf_ram.memory\[273\]\[1\] _05181_ _05183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_204_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_196_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11432__A1 _04817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14350_ _00204_ net3 mod.u_cpu.rf_ram.memory\[512\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_195_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_196_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13301_ _06383_ _06362_ _06375_ _06396_ _06398_ _06399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_168_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10513_ _04452_ _04469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_11_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14281_ _00135_ net3 mod.u_cpu.rf_ram.memory\[547\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11493_ _05114_ mod.u_cpu.rf_ram.memory\[284\]\[0\] _05136_ _05137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_137_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13232_ _06338_ _06339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_10444_ _04421_ _00326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_108_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07939__A1 _02245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13468__I _06512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15331__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13163_ _06204_ _06273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_10375_ _04365_ mod.u_cpu.rf_ram.memory\[462\]\[0\] _04374_ _04375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08600__A2 mod.u_cpu.rf_ram.memory\[262\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10794__I0 _04641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07466__I _01744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12114_ _05558_ _00859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_174_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_112_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13094_ _06230_ mod.u_cpu.rf_ram.memory\[59\]\[0\] _06231_ _06232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_152_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12045_ _05488_ _05512_ _05513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_215_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07167__A2 _01471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15481__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08364__A1 _02638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12160__A2 _05589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_266_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_265_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_238_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_226_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11716__I _05249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10620__I _04541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_207_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_207_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13996_ _06957_ _06959_ _01340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_19_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12947_ _03500_ mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat\[0\] _06124_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_3171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_3182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13931__I _05801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_206_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_234_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_222_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_244_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12878_ _06075_ _01106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_178_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14617_ _00471_ net3 mod.u_cpu.rf_ram.memory\[37\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_92_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11829_ _05328_ _05364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_53_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11451__I _05105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15597_ _01368_ net3 mod.u_cpu.rf_ram.memory\[245\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13412__A2 _06011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_187_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_222_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_144_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_187_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14548_ _00402_ net3 mod.u_cpu.rf_ram.memory\[413\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_187_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09092__A2 _03392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14429__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11974__A2 _04108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_174_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14479_ _00333_ net3 mod.u_cpu.rf_ram.memory\[448\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_146_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_31_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_127_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12774__I1 _06005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_255_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14579__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_170_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08971_ mod.u_cpu.cpu.bufreg2.i_cnt_done _03272_ _03273_ _03275_ _03276_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_102_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_229_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07922_ _01719_ _02230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_9_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07158__A2 _01465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09591__I _03804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_256_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07853_ _01646_ _02161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_217_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14002__I _06963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_244_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07784_ _02091_ _02092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_09523_ _03271_ _03715_ _03705_ _01461_ _03747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_25_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_65_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11562__S _05181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13651__A2 _06662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_213_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09454_ _03255_ _03681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_197_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15204__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10465__A2 _04132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_266_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_197_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_240_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_101_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08405_ mod.u_cpu.rf_ram.memory\[440\]\[1\] mod.u_cpu.rf_ram.memory\[441\]\[1\] mod.u_cpu.rf_ram.memory\[442\]\[1\]
+ mod.u_cpu.rf_ram.memory\[443\]\[1\] _02711_ _01703_ _02712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_52_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09385_ _03563_ _03623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_24_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13403__A2 _06403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_212_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11414__A1 _04804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08336_ _02631_ _02634_ _02642_ _01587_ _02643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_177_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_193_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07713__S0 _02020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__15354__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08267_ _02546_ mod.u_cpu.rf_ram.memory\[540\]\[0\] _02574_ _02575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_193_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09766__I _03697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07218_ _01517_ mod.u_cpu.rf_ram.memory\[454\]\[0\] _01522_ _01525_ _01526_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_118_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08198_ _02449_ _02496_ _02504_ _02505_ _02506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_134_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07149_ _01457_ _01458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_195_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10160_ mod.u_cpu.cpu.immdec.imm11_7\[4\] _04222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_134_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_120_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_266_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_248_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10091_ _04136_ _04173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08346__A1 _01592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_247_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08897__A2 _03196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_75_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13850_ _06472_ _06443_ _06466_ _06845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_210_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_263_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_216_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12801_ _03985_ _06011_ _06024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_28_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_262_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_13781_ _06381_ _06372_ _06781_ _06782_ _06432_ _06783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_10993_ _04792_ _04788_ _04793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_216_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15520_ _01291_ net3 mod.u_cpu.cpu.immdec.imm31 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_128_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12732_ _03932_ _05978_ _05979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_216_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_203_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_245_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07321__A2 _01621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_204_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15451_ _01225_ net3 mod.u_cpu.cpu.ctrl.o_ibus_adr\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_71_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_230_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10088__S _04169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12663_ _05923_ mod.u_cpu.rf_ram.memory\[144\]\[1\] _05931_ _05933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_208_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14402_ _00256_ net3 mod.u_cpu.rf_ram.memory\[486\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11614_ _05208_ mod.u_cpu.rf_ram.memory\[264\]\[1\] _05215_ _05217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_54_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15382_ _01157_ net3 mod.u_cpu.rf_ram.memory\[106\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_169_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12594_ _05886_ _05887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_211_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14333_ _00187_ net3 mod.u_cpu.rf_ram.memory\[521\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11545_ _05124_ _05171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_129_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08821__A2 mod.u_cpu.rf_ram.memory\[30\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09676__I _03871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14721__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11476_ _05118_ _05124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_14264_ _00118_ net3 mod.u_cpu.rf_ram.memory\[555\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_144_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12905__A1 _05657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13215_ _06286_ _06287_ _06322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_143_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10427_ _04344_ _04410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_100_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10767__I0 _04637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14195_ _07076_ _07094_ _01404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__07196__I _01503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08585__A1 _01992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_252_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13146_ mod.u_arbiter.i_wb_cpu_rdt\[24\] mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat\[8\]
+ _06263_ _06264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_152_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10358_ _04344_ _04363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_124_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14871__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_151_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13077_ _06220_ _01160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_183_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10289_ _04298_ mod.u_cpu.rf_ram.memory\[476\]\[0\] _04316_ _04317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__13330__A1 _06316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_238_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_12028_ _05502_ _00829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08888__A2 _03187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_211_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_266_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15227__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10695__A2 _04575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_226_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14130__I0 _07041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07560__A2 mod.u_cpu.rf_ram.memory\[382\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_253_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_207_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_202_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13979_ _06910_ _06947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_47_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_18_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_222_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14251__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15377__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_222_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09170_ mod.u_arbiter.i_wb_cpu_rdt\[13\] mod.u_arbiter.i_wb_cpu_dbus_dat\[10\] _03452_
+ _03455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_203_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08121_ _02329_ mod.u_cpu.rf_ram.memory\[36\]\[0\] _02428_ _02429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08112__I1 mod.u_cpu.rf_ram.memory\[53\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08052_ _02356_ mod.u_cpu.rf_ram.memory\[70\]\[0\] _02358_ _02359_ _02360_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_107_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_128_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10758__I0 _04626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08576__A1 _01979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_153_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10383__A1 _04377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12740__I _05937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08954_ _03258_ _03259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_130_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_257_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07905_ _02211_ mod.u_cpu.rf_ram.memory\[210\]\[0\] _02212_ _02213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_4619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08885_ _02500_ _03191_ _03192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_116_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_229_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13872__A2 mod.u_arbiter.i_wb_cpu_rdt\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3907 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10260__I _04250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3918 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07836_ _02124_ _02128_ _02142_ _02143_ _02144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_99_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_245_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3929 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07767_ mod.u_cpu.rf_ram.memory\[156\]\[0\] mod.u_cpu.rf_ram.memory\[157\]\[0\] mod.u_cpu.rf_ram.memory\[158\]\[0\]
+ mod.u_cpu.rf_ram.memory\[159\]\[0\] _01925_ _02071_ _02075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_112_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_213_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_266_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09506_ _01462_ mod.u_cpu.rf_ram_if.wdata1_r\[1\] _03731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_37_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07698_ _01997_ _02001_ _02004_ _02005_ _02006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_77_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__07303__A2 mod.u_cpu.rf_ram.memory\[508\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_198_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_227_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_197_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09437_ _03289_ _03667_ _03668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_212_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__07502__C _01783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_213_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__14744__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12435__I0 mod.u_cpu.rf_ram.memory\[173\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09368_ _03386_ mod.u_scanchain_local.module_data_in\[59\] _03401_ mod.u_arbiter.i_wb_cpu_dbus_adr\[22\]
+ _03609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_40_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_166_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_205_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08319_ _02198_ mod.u_cpu.rf_ram.memory\[470\]\[1\] _02625_ _01751_ _02626_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_177_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09299_ _03535_ mod.u_scanchain_local.module_data_in\[48\] _03536_ mod.u_arbiter.i_wb_cpu_dbus_adr\[11\]
+ _03551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__08803__A2 _03109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14188__I0 _03699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_197_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11330_ _05007_ mod.u_cpu.rf_ram.memory\[310\]\[0\] _05025_ _05026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_20_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_165_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14894__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11261_ _04977_ _00587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_181_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08567__A1 _01848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10212_ _04245_ mod.u_cpu.rf_ram.memory\[487\]\[1\] _04259_ _04261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_106_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13000_ _06113_ _06166_ _06170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_140_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11410__I1 _04954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11192_ _03909_ _04930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_84_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_97_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10374__A1 _04218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10143_ _04193_ mod.u_cpu.rf_ram.memory\[496\]\[0\] _04210_ _04211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08319__A1 _02198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13312__A1 _06401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_251_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14951_ _00805_ net3 mod.u_cpu.rf_ram.memory\[218\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10074_ _04157_ mod.u_cpu.rf_ram.memory\[506\]\[1\] _04159_ _04161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_94_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_212_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__13863__A2 _06836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13902_ _03359_ _06422_ _06693_ _06463_ _06699_ _06135_ _01320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai222_1
XFILLER_134_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_208_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14882_ _00736_ net3 mod.u_cpu.rf_ram.memory\[242\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_63_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14274__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13833_ _06764_ _06829_ _06830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_235_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12298__S _05683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_204_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_216_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_262_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13764_ mod.u_cpu.cpu.immdec.imm19_12_20\[8\] _06767_ _06709_ _06768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_10976_ _04414_ _04781_ _04782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_204_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07925__S0 _02151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_16_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_15503_ _01274_ net3 mod.u_arbiter.i_wb_cpu_dbus_adr\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_189_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08508__C _01687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12715_ _03918_ _05940_ _05968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_231_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_204_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13695_ _05787_ _06704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_30_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_188_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15434_ _01209_ net3 mod.u_cpu.cpu.immdec.imm11_7\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12646_ _05922_ _01027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_178_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14040__A2 _06989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15365_ _01140_ net3 mod.u_cpu.rf_ram.memory\[10\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_157_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12577_ _05428_ _05374_ _05876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10988__I0 _04774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_200_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14316_ _00170_ net3 mod.u_cpu.rf_ram.memory\[52\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_144_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11528_ _04741_ _05149_ _05160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_184_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15296_ _00056_ net4 mod.u_scanchain_local.module_data_in\[53\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_183_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14247_ _00101_ net3 mod.u_cpu.rf_ram.memory\[564\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11459_ _05112_ _00650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_256_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12354__A2 _05721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11401__I1 mod.u_cpu.rf_ram.memory\[2\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14178_ _07057_ mod.u_cpu.rf_ram.memory\[8\]\[0\] _07083_ _07084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_139_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13129_ _06254_ _01178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07654__I _01752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12106__A2 _05553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_239_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14617__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11165__I0 _04896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08405__S1 _01703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_113_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_152_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08670_ _02759_ _02973_ _02976_ _01872_ _02977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_94_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08686__S _01545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_227_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08730__A1 _02043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14103__I0 _07028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07621_ _01686_ _01929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_66_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_214_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11617__A1 _05133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07552_ _01858_ _01859_ _01860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__14767__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_207_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_228_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_222_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07483_ _01445_ _01791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_222_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09222_ _03435_ mod.u_scanchain_local.module_data_in\[37\] _03485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_210_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10840__A2 _04687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_188_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09153_ mod.u_arbiter.i_wb_cpu_dbus_dat\[4\] _03444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_147_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13090__I0 _06217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08104_ mod.u_cpu.rf_ram.memory\[23\]\[0\] _02412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__08797__A1 _02348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09084_ _03384_ _03385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_108_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11640__I1 mod.u_cpu.rf_ram.memory\[260\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08035_ _01662_ _02342_ _02343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_190_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12470__I _05709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09986_ _04013_ _03851_ _04100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_5117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_118_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14297__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_233_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08937_ _03234_ _03243_ _02520_ _03244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_4416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15542__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_218_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08868_ _02455_ _03171_ _03174_ _02555_ _03175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_3726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08721__A1 _02591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_217_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07819_ _02126_ _02127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_3759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08799_ mod.u_cpu.rf_ram.memory\[69\]\[1\] _03106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_38_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_244_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12656__I0 _05918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10830_ _04681_ _00452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_38_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_260_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_198_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_198_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10761_ _04622_ mod.u_cpu.rf_ram.memory\[3\]\[0\] _04634_ _04635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_12_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12500_ _05822_ mod.u_cpu.rf_ram.memory\[459\]\[1\] _05824_ _05826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_164_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_198_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13480_ _03598_ _06545_ _06546_ _03602_ _06547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_10692_ _04589_ _00406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_199_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_197_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_240_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_201_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12431_ _05773_ _00961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_225_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_194_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07739__I _02026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_194_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13781__A1 _06381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15150_ _01003_ net3 mod.u_cpu.rf_ram.memory\[15\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12362_ _05713_ mod.u_cpu.rf_ram.memory\[180\]\[0\] _05727_ _05728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_165_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14101_ _07021_ mod.u_cpu.rf_ram.memory\[110\]\[0\] _07033_ _07034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_11313_ _04951_ _05014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10165__I _04226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15081_ _00935_ net3 mod.u_cpu.rf_ram.memory\[181\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12293_ _05679_ mod.u_cpu.rf_ram.memory\[188\]\[0\] _05680_ _05681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_107_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15072__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11244_ _04965_ _04945_ _04966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_14032_ mod.u_arbiter.i_wb_cpu_dbus_dat\[22\] _06978_ _06986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_107_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11395__I0 _05069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_122_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11175_ _04775_ _04906_ _04919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_136_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07474__I _01700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10126_ _04177_ _04199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_122_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_95_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_209_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07407__C _01714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_248_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13836__A2 _06774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_209_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14934_ _00788_ net3 mod.u_cpu.rf_ram.memory\[225\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10057_ _04150_ _00210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11698__I1 mod.u_cpu.rf_ram.memory\[254\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4950 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_212_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_264_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08712__A1 _03017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4961 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07366__I2 mod.u_cpu.rf_ram.memory\[390\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4972 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_180_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4983 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14865_ _00719_ net3 mod.u_cpu.rf_ram.memory\[250\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_169_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4994 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_90_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13816_ mod.u_arbiter.i_wb_cpu_rdt\[28\] mod.u_arbiter.i_wb_cpu_rdt\[12\] _03510_
+ _06815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_63_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_263_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14796_ _00650_ net3 mod.u_cpu.rf_ram.memory\[28\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09268__A2 _03521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_204_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13747_ _06752_ _01298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__12272__A1 _03755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10959_ _04769_ _00493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_250_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_232_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_204_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10822__A2 _03951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_177_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13678_ _06421_ _06688_ _06689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_148_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15417_ _01192_ net3 mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_12629_ _05907_ mod.u_cpu.rf_ram.memory\[150\]\[1\] _05909_ _05911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_223_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08779__A1 _01688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07649__I _01919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15415__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15348_ _01123_ net3 mod.u_cpu.rf_ram.memory\[379\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_184_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09440__A2 _03331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_258_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_145_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15279_ _00037_ net4 mod.u_scanchain_local.module_data_in\[36\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_144_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_172_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09864__I _03762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_217_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_63_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08701__C _01669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15565__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09840_ _04000_ _00143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_99_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10803__I _04621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10889__A2 _04722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09771_ _03947_ _00127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_100_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13827__A2 _06324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_230_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08722_ _03016_ _03019_ _02074_ _03028_ _03029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_227_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08653_ _02135_ mod.u_cpu.rf_ram.memory\[166\]\[1\] _02959_ _02139_ _02960_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_254_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_227_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_227_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_226_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07604_ _01848_ _01889_ _01911_ _01912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__14010__I _06909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_199_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08584_ _01997_ _02887_ _02890_ _02005_ _02891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_81_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_242_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09104__I _03403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_223_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07535_ _01825_ _01843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_228_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_179_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_263_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07466_ _01744_ _01774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_168_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_210_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09205_ _03475_ _00031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_241_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07397_ _01704_ _01705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_249_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_195_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15095__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07559__I _01503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_210_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09136_ _03430_ _03431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_159_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09067_ _03353_ _03369_ _03370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_136_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_191_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09774__I _03949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_191_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08018_ mod.u_cpu.rf_ram.memory\[117\]\[0\] _02326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__07993__A2 mod.u_cpu.rf_ram.memory\[108\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_239_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08617__S1 _02043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07508__B _01738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07294__I _01492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14932__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07227__C _01534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09969_ _04073_ mod.u_cpu.rf_ram.memory\[522\]\[0\] _04088_ _04089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_249_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13818__A2 _06816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_218_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_134_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_170_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12877__I0 _06073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12980_ mod.u_cpu.cpu.decode.op22 _03343_ _06151_ _06154_ _06155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XTAP_4246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13294__A3 _06391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09215__S _03479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_218_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11931_ _03698_ _05437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_3534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09442__C _03672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_175_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10501__A1 _04322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14650_ _00504_ net3 mod.u_cpu.rf_ram.memory\[362\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12629__I0 _05907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11862_ _05387_ _05388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_233_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13601_ mod.u_cpu.rf_ram.memory\[329\]\[0\] _03899_ _06621_ _06622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_26_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_261_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12254__A1 _05408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_207_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10813_ _04663_ mod.u_cpu.rf_ram.memory\[391\]\[0\] _04670_ _04671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_2877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14581_ _00435_ net3 mod.u_cpu.rf_ram.memory\[397\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11793_ _05340_ _00756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11301__I0 _04999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2899 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10104__I1 mod.u_cpu.rf_ram.memory\[502\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_232_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14312__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_198_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15438__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13532_ _03292_ _06583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_10744_ _04201_ _04623_ _04624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_198_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13463_ _06535_ _01231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_201_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10675_ _04496_ _04578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_142_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15202_ _01055_ net3 mod.u_cpu.rf_ram.memory\[78\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09885__S _04030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13754__A1 _06432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12414_ _05762_ _00955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_167_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13394_ _06485_ _06488_ _06489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_182_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08076__I3 mod.u_cpu.rf_ram.memory\[7\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14462__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15133_ _00986_ net3 mod.u_cpu.rf_ram.memory\[166\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__15588__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_182_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12345_ _05711_ mod.u_cpu.rf_ram.memory\[182\]\[1\] _05714_ _05716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_181_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09684__I _03809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13506__A1 _06142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07984__A2 _02282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15064_ _00918_ net3 mod.u_cpu.rf_ram.memory\[187\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_142_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12276_ _05662_ mod.u_cpu.rf_ram.memory\[191\]\[0\] _05669_ _05670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_107_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08608__S1 _02067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11719__I _05221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14015_ mod.u_arbiter.i_wb_cpu_rdt\[16\] _06964_ _06971_ mod.u_arbiter.i_wb_cpu_dbus_dat\[16\]
+ _06974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_11227_ _04953_ _00577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_136_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_253_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08933__A1 _02551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11158_ _04901_ mod.u_cpu.rf_ram.memory\[337\]\[0\] _04907_ _04908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_136_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_209_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_249_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10109_ _04186_ _04185_ _04187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_11089_ _04843_ mod.u_cpu.rf_ram.memory\[348\]\[0\] _04860_ _04861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_67_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09489__A2 _03374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14917_ _00771_ net3 mod.u_cpu.rf_ram.memory\[228\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_236_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13690__B1 _06699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_224_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_209_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_208_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14848_ _00702_ net3 mod.u_cpu.rf_ram.memory\[263\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_63_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11048__A2 _04822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_210_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14779_ _00633_ net3 mod.u_cpu.rf_ram.memory\[298\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__13293__I0 mod.u_arbiter.i_wb_cpu_rdt\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_182_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08839__I2 _03144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_251_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09859__I _03809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07320_ _01572_ _01624_ _01627_ _01584_ _01628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__13993__A1 mod.u_arbiter.i_wb_cpu_dbus_dat\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12796__A2 _03905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_177_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_260_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_108_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07251_ _01556_ mod.u_cpu.rf_ram.memory\[476\]\[0\] _01558_ _01559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_220_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14805__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13045__I0 _06199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_220_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07600__C _01882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_192_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07379__I _01686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07182_ mod.u_cpu.raddr\[2\] _01490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_191_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_121_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08847__S1 _01732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_258_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08712__B _01870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14955__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14170__A1 _06047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12020__I1 mod.u_cpu.rf_ram.memory\[214\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14005__I _06942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08924__A1 _02534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09823_ _03767_ _03986_ _03987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_99_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10582__I1 mod.u_cpu.rf_ram.memory\[42\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11565__S _05184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_189_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09754_ _03902_ _03933_ _03934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07842__I _01741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09024__S1 mod.u_cpu.cpu.bufreg.lsb\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08705_ mod.u_cpu.rf_ram.memory\[238\]\[1\] mod.u_cpu.rf_ram.memory\[239\]\[1\] _01807_
+ _03012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_104_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11287__A2 _04996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_261_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09685_ _03822_ _03879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_54_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_255_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08152__A2 mod.u_cpu.rf_ram.memory\[548\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14335__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_227_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08636_ _01836_ _02940_ _02942_ _02943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_243_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08567_ _01848_ _02854_ _02873_ _02874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_120_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_214_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_154_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_230_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08535__S0 _01753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10098__I0 _04178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_211_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07518_ _01825_ _01826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_165_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08498_ _01875_ mod.u_cpu.rf_ram.memory\[334\]\[1\] _02804_ _02453_ _02805_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_126_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__14485__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07663__A1 _01697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_195_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07449_ _01515_ _01757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_168_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_210_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13736__A1 _06726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_182_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10460_ _04290_ _04309_ _04432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13736__B2 _06442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09404__A2 _03615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08838__S1 _02388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_182_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09119_ _03416_ _03392_ _03417_ _03418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_10391_ _04386_ _00308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12923__I _06017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_237_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_191_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12130_ _05559_ mod.u_cpu.rf_ram.memory\[208\]\[0\] _05569_ _05570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_159_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12061_ _05518_ mod.u_cpu.rf_ram.memory\[62\]\[1\] _05522_ _05524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_78_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08915__A1 _02550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11012_ _04797_ mod.u_cpu.rf_ram.memory\[360\]\[1\] _04805_ _04807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09963__I0 _04073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15110__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10573__I1 mod.u_cpu.rf_ram.memory\[430\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08391__A2 mod.u_cpu.rf_ram.memory\[422\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4010 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4021 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4032 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_253_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4043 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4054 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4065 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12963_ _06139_ _06140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12475__A1 _05759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_218_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_4076 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4087 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4098 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14702_ _00556_ net3 mod.u_cpu.rf_ram.memory\[336\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_46_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11914_ _05425_ _00792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15260__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12894_ _06085_ _01112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14633_ _00487_ net3 mod.u_cpu.rf_ram.memory\[371\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__14828__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11845_ _05376_ _00772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1940 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_220_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1951 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_233_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1962 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_207_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14564_ _00418_ net3 mod.u_cpu.rf_ram.memory\[405\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1973 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11776_ _05328_ _05329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_207_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1984 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1995 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_198_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_158_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13515_ _03693_ _06568_ _06569_ _06570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_159_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10727_ _01725_ _04610_ _04612_ _00418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_202_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14495_ _00349_ net3 mod.u_cpu.rf_ram.memory\[440\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_186_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14978__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13446_ _06510_ _06525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_70_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10658_ _04557_ mod.u_cpu.rf_ram.memory\[416\]\[0\] _04565_ _04566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__11589__I0 _05199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_127_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13377_ _06471_ _06464_ _06458_ _06395_ _06472_ _06473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_103_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10589_ _04238_ _04507_ _04519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_155_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07957__A2 _02257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15116_ _00969_ net3 mod.u_cpu.rf_ram.memory\[519\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_127_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12328_ _05283_ _05703_ _05704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_181_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10961__A1 _04746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15047_ _00901_ net3 mod.u_cpu.rf_ram.memory\[196\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_64_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12259_ _03979_ _05657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_69_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07709__A2 mod.u_cpu.rf_ram.memory\[262\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_214_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12702__A2 _04643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10713__A1 _04172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11761__I0 _05304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14358__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07662__I _01701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15603__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_243_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_237_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11513__I0 _05144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xtiny_user_project_170 wbs_dat_o[20] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_225_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xtiny_user_project_181 wbs_dat_o[31] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__08134__A2 _02438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_184_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_209_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09470_ _03695_ _03696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_52_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__14207__A2 _05210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_221_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08421_ _02244_ _02727_ _02728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_97_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07893__A1 _02198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_212_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_264_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_196_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08352_ _02656_ _02657_ _02658_ _02067_ _02659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_189_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07303_ _01607_ mod.u_cpu.rf_ram.memory\[508\]\[0\] _01610_ _01611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07645__A1 _01938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08283_ _02561_ _02586_ _02589_ _02080_ _02590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_20_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07234_ mod.u_cpu.rf_ram.memory\[461\]\[0\] _01542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_146_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_192_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13194__A2 _06300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07165_ _01472_ _01473_ _01474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_146_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10252__I0 _04288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08070__A1 _02365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11359__I _04959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15133__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_160_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_161_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09806_ _03973_ _03974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_115_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15283__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07998_ _01569_ _02306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_235_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_228_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09737_ _03916_ mod.u_cpu.rf_ram.memory\[554\]\[0\] _03920_ _03921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_101_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07505__C _01812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11094__I _04802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09668_ _03865_ _03866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_27_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_215_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08619_ mod.u_cpu.rf_ram.memory\[152\]\[1\] mod.u_cpu.rf_ram.memory\[153\]\[1\] mod.u_cpu.rf_ram.memory\[154\]\[1\]
+ mod.u_cpu.rf_ram.memory\[155\]\[1\] _02066_ _02067_ _02926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__13406__B1 _06498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09599_ _03812_ _00090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_202_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_215_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11630_ _04817_ _05227_ _05228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_39_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_208_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08336__C _01587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_196_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07636__A1 _01791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11561_ _05182_ _00682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_129_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07240__C _01525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13709__A1 _06380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13300_ _06397_ _06398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_10_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10512_ _04468_ _00347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10491__I0 _04453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14280_ _00134_ net3 mod.u_cpu.rf_ram.memory\[547\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_155_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11492_ _04859_ _05125_ _05136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_109_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_196_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13231_ _06337_ _06338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_137_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10443_ _04400_ mod.u_cpu.rf_ram.memory\[451\]\[0\] _04420_ _04421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_6_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12232__I1 _05617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_170_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08352__B _02658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_13162_ _06272_ _01193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_174_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_136_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10374_ _04218_ _04373_ _04374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_108_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_163_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12113_ _05550_ mod.u_cpu.rf_ram.memory\[68\]\[1\] _05556_ _05558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_124_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10173__I _03904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13093_ _05888_ _03878_ _06231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_123_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__14500__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15626__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12044_ _05164_ _05433_ _05512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07247__S0 _01540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_266_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_104_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07167__A3 _01475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08364__A2 mod.u_cpu.rf_ram.memory\[484\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_211_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_225_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12448__A1 mod.u_arbiter.i_wb_cpu_ibus_adr\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13995_ mod.u_arbiter.i_wb_cpu_rdt\[11\] _06952_ _06958_ mod.u_arbiter.i_wb_cpu_dbus_dat\[11\]
+ _06959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__14650__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_219_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_234_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_234_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_207_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12946_ mod.u_arbiter.i_wb_cpu_rdt\[0\] _06123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XTAP_3161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_206_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07875__A1 _02179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_209_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_12877_ _06073_ mod.u_cpu.rf_ram.memory\[246\]\[0\] _06074_ _06075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_61_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_234_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_221_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08527__B _02040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15006__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14616_ _00470_ net3 mod.u_cpu.rf_ram.memory\[37\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_33_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11828_ _02430_ _05362_ _05363_ _00768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_15596_ _01367_ net3 mod.u_cpu.rf_ram.memory\[245\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__14070__B1 _06919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_261_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08246__C _02515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14547_ _00401_ net3 mod.u_cpu.rf_ram.memory\[414\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11759_ _05265_ _05316_ _05317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_18_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12620__A1 _03879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_186_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_197_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_146_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14478_ _00332_ net3 mod.u_cpu.rf_ram.memory\[448\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_186_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__15156__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13429_ _06515_ _01217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__13420__I0 _06354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11187__A1 _04784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_220_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08052__A1 _02356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08970_ mod.u_cpu.cpu.bufreg2.i_cnt_done mod.u_cpu.cpu.immdec.imm31 _03274_ _03275_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_130_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07921_ _02120_ _02214_ _02219_ _02224_ _02228_ _02229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_142_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07852_ _02156_ mod.u_cpu.rf_ram.memory\[196\]\[0\] _02159_ _02160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07392__I _01497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10162__A2 _03753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput1 io_in[10] net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_84_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07783_ _01671_ _02091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_72_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09522_ _01850_ _03703_ _03746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_83_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_225_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_225_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_213_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09453_ _03395_ _03679_ _03680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_80_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_149_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_08404_ _01518_ _02711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_197_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09384_ _03613_ _03622_ _00066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_101_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_178_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08335_ _02597_ _02637_ _02641_ _01651_ _02642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__11414__A2 _05058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07713__S1 _01995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08266_ _02472_ _02573_ _02574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_192_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13569__I _03692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_197_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07217_ _01524_ _01525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_119_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_193_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_257_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_197_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08197_ _02122_ _02505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_180_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07567__I _01825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_238_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14523__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07148_ _01450_ _01456_ _01457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_69_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10925__A1 _04746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10776__I1 _04396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_133_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09918__I0 _04054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10090_ _03821_ _04172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_160_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14673__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10721__I _04578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_248_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_207_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_262_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_216_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12800_ _06023_ _01080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__15029__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13780_ _06494_ _06324_ _06380_ _06782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_90_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11102__A1 _04868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10992_ _03917_ _04792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_55_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12731_ _05919_ _05978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_231_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07857__A1 _02161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_255_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_231_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12850__A1 _02505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_204_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_203_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15450_ _01224_ net3 mod.u_cpu.cpu.ctrl.o_ibus_adr\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12662_ _05932_ _01033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_187_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_231_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15179__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14401_ _00255_ net3 mod.u_cpu.rf_ram.memory\[487\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_231_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11613_ _05216_ _00700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12602__A1 _03796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10168__I _03898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15381_ _01156_ net3 mod.u_cpu.rf_ram.memory\[106\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_180_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12593_ _05694_ _05886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_129_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14332_ _00186_ net3 mod.u_cpu.rf_ram.memory\[521\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11544_ _05170_ _00677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_156_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08282__A1 _02560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_204_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__13479__I _06539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_184_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14263_ _00117_ net3 mod.u_cpu.rf_ram.memory\[556\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11475_ _05123_ _00655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_167_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07477__I _01765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13214_ _06320_ _06321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_167_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10426_ _04409_ _00320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12905__A2 _06092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14194_ _07067_ _03389_ _03674_ _07093_ _07094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__11964__I0 _05442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10767__I1 mod.u_cpu.rf_ram.memory\[398\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08585__A2 _02884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_174_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_13145_ _06252_ _06263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_10357_ _04362_ _00298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_112_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_140_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_174_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13076_ mod.u_cpu.rf_ram.memory\[105\]\[0\] _05971_ _06219_ _06220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_215_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10288_ _04315_ _04303_ _04316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_78_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12027_ _05501_ mod.u_cpu.rf_ram.memory\[58\]\[1\] _05499_ _05502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__13330__A2 _06426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_266_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07426__B _01733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_266_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_265_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_254_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_250_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_226_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_219_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13978_ mod.u_arbiter.i_wb_cpu_dbus_dat\[8\] _06943_ _06946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_47_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_234_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_207_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12929_ _06107_ mod.u_cpu.rf_ram.memory\[369\]\[0\] _06108_ _06109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__11462__I _05045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_179_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_210_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_107_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_222_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10078__I _04142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_194_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15579_ _01350_ net3 mod.u_arbiter.i_wb_cpu_dbus_dat\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_187_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_175_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08120_ _02406_ _02427_ _02428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__14546__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08273__A1 _02542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08051_ _01820_ _02359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_135_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_257_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_174_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_190_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07387__I _01491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_179_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10207__I0 _04245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08025__A1 _02325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_192_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__14696__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08576__A2 _02875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10383__A2 _04380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_170_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_248_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_170_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08953_ mod.u_cpu.cpu.mem_bytecnt\[0\] mod.u_cpu.cpu.state.o_cnt\[2\] mod.u_cpu.cpu.mem_bytecnt\[1\]
+ _03258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_9_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07904_ _01701_ _02212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10541__I _04442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08884_ mod.u_cpu.rf_ram.memory\[575\]\[1\] _03191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_111_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12380__I0 _05731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_217_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3908 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07835_ _01533_ _02143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3919 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_244_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11573__S _05188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_186_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07766_ _01890_ _02074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08946__I _01421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12132__I0 _05566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_260_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09828__A2 _03818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_225_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09505_ _03730_ _00078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07839__A1 _02103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_213_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_198_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15321__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_198_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07697_ _01491_ _02005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_80_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08500__A2 _02799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_240_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09436_ mod.u_cpu.cpu.state.init_done _01434_ _03667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__09978__S _04093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_52_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_25_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_198_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_80_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_201_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09367_ _03605_ _03606_ _03608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__12435__I1 _05765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_205_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_200_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08318_ _02115_ _02624_ _02625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_162_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15471__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09298_ _03547_ _03548_ _03549_ _03550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_193_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13299__I _06328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10071__A1 _03797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08249_ _02542_ _02544_ _02556_ _02491_ _02557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_126_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_193_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07297__I _01604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_180_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11260_ _04976_ mod.u_cpu.rf_ram.memory\[321\]\[1\] _04974_ _04977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12899__A1 _03985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_134_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10211_ _01625_ _04259_ _04260_ _00254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_137_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11191_ _04929_ _00565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_107_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11571__A1 _05133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_234_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10142_ _04209_ _04202_ _04210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08319__A2 mod.u_cpu.rf_ram.memory\[470\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14950_ _00804_ net3 mod.u_cpu.rf_ram.memory\[218\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10073_ _04160_ _00216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_212_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__11323__A1 _05019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_247_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_236_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_13901_ _03306_ _06881_ _06689_ _01319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_14881_ _00735_ net3 mod.u_cpu.rf_ram.memory\[243\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_169_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14419__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_263_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13832_ _05790_ _03670_ _03679_ _06829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_75_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12123__I0 _05559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_210_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13763_ _06761_ _06763_ _06765_ _06766_ _06767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_10975_ _04377_ _04780_ _04781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_216_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_44_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_245_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__07925__S1 _02172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12714_ _05967_ _01050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__14569__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15502_ _01273_ net3 mod.u_arbiter.i_wb_cpu_dbus_adr\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_13694_ _06703_ _01294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_71_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15433_ _01208_ net3 mod.u_cpu.cpu.immdec.imm11_7\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_176_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12645_ _05918_ mod.u_cpu.rf_ram.memory\[147\]\[0\] _05921_ _05922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__13623__I0 _06581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_169_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_15364_ _01139_ net3 mod.u_cpu.rf_ram.memory\[85\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_157_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12576_ _05875_ _01004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_30_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_200_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08524__C _01867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14315_ _00169_ net3 mod.u_cpu.rf_ram.memory\[530\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11527_ _05143_ _05159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_183_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15295_ _00055_ net4 mod.u_scanchain_local.module_data_in\[52\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_171_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14246_ _00100_ net3 mod.u_cpu.rf_ram.memory\[564\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_183_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08007__A1 _02297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11458_ _05096_ mod.u_cpu.rf_ram.memory\[28\]\[0\] _05111_ _05112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_125_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13000__A1 _06113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13937__I _05792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10409_ _04398_ _00314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_14177_ _06181_ _03933_ _07083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11389_ mod.u_cpu.rf_ram.memory\[301\]\[1\] _05065_ _05063_ _05066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_113_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_259_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_13128_ mod.u_arbiter.i_wb_cpu_rdt\[16\] mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat\[0\]
+ _06253_ _06254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_152_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_140_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09507__A1 _01462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10361__I _04347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13059_ _04107_ _05589_ _06209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_140_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_152_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_61_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_39_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12362__I0 _05713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_227_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_16_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15344__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_227_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_226_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07620_ _01925_ mod.u_cpu.rf_ram.memory\[318\]\[0\] _01927_ _01783_ _01928_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_253_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_242_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07670__I _01832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_263_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12288__I _05634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07551_ mod.u_cpu.rf_ram.memory\[381\]\[0\] _01859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__12814__A1 _06032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11192__I _03909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_222_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08494__A1 _01729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15494__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07482_ _01740_ _01769_ _01789_ _01790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_195_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09221_ _03483_ _03435_ _03484_ _00038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_107_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_188_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10428__I0 _04410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09152_ _03443_ _00077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08246__A1 _02550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_175_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_238_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08103_ _01778_ _02411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08434__C _01658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08797__A2 _03103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09083_ net2 _03384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_190_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_200_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08034_ mod.u_cpu.rf_ram.memory\[88\]\[0\] mod.u_cpu.rf_ram.memory\[89\]\[0\] mod.u_cpu.rf_ram.memory\[90\]\[0\]
+ mod.u_cpu.rf_ram.memory\[91\]\[0\] _01673_ _01666_ _02342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_174_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_192_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_192_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08450__B _01483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_89_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_35 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_235_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_249_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_235_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09985_ _04099_ _00189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_5118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10271__I _04302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08936_ _02542_ _03235_ _03242_ _02518_ _03243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_88_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_229_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_218_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_218_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08867_ _02461_ mod.u_cpu.rf_ram.memory\[550\]\[1\] _03173_ _02578_ _03174_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_111_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_123_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_245_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08721__A2 _03020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07818_ _01568_ _02126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08798_ mod.u_cpu.rf_ram.memory\[64\]\[1\] mod.u_cpu.rf_ram.memory\[65\]\[1\] mod.u_cpu.rf_ram.memory\[66\]\[1\]
+ mod.u_cpu.rf_ram.memory\[67\]\[1\] _01561_ _01714_ _03105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__14711__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_226_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_26_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07749_ _01487_ _02057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_226_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_198_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_241_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10760_ _04196_ _03969_ _04634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07288__A2 mod.u_cpu.rf_ram.memory\[500\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_242_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09419_ _03439_ mod.u_scanchain_local.module_data_in\[66\] _03653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_158_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14861__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10691_ _04584_ mod.u_cpu.rf_ram.memory\[411\]\[0\] _04588_ _04589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_201_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12430_ _05761_ mod.u_cpu.rf_ram.memory\[439\]\[1\] _05771_ _05773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_90_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_200_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13230__A1 _06137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_201_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11092__I0 _04862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08344__C _01651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13781__A2 _06372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12361_ _05535_ _05726_ _05727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_120_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_218_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_148_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15217__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14100_ _03885_ _07014_ _07033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11312_ _05013_ _00602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_154_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15080_ _00934_ net3 mod.u_cpu.rf_ram.memory\[181\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_181_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_148_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12292_ _05443_ _05668_ _05680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_180_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_153_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14031_ _06984_ _06985_ _01349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_153_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11243_ _03967_ _04965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08096__S0 _02403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11395__I1 mod.u_cpu.rf_ram.memory\[300\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11174_ _04882_ _04918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_136_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14241__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15367__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11277__I _04988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10125_ _04198_ _00230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11147__I1 _04819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_236_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14933_ _00787_ net3 mod.u_cpu.rf_ram.memory\[226\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10056_ _04148_ mod.u_cpu.rf_ram.memory\[50\]\[0\] _04149_ _04150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_208_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4940 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4951 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4962 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_180_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08712__A2 _03018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4973 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12102__S _05547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13049__A1 _02373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14391__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_235_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_224_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14864_ _00718_ net3 mod.u_cpu.rf_ram.memory\[250\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_4984 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_224_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4995 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13815_ _06431_ _06814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_14795_ _00649_ net3 mod.u_cpu.rf_ram.memory\[290\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_169_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_204_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_204_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10658__I0 _04557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13746_ mod.u_cpu.cpu.immdec.imm19_12_20\[6\] _06658_ _06749_ _06751_ _06752_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_16_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__12272__A2 _05371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10958_ _04756_ mod.u_cpu.rf_ram.memory\[368\]\[1\] _04767_ _04769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_204_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_231_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_188_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_177_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13677_ _06451_ _06685_ _06687_ _06688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__12836__I _06046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10889_ _04414_ _04722_ _04723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_108_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_15416_ _01191_ net3 mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12628_ _05910_ _01021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08228__A1 _02534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_176_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_169_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_185_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10035__A1 mod.u_cpu.cpu.immdec.imm11_7\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_185_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11083__I0 _04843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15347_ _01122_ net3 mod.u_cpu.rf_ram.memory\[379\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_184_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12559_ _05855_ mod.u_cpu.rf_ram.memory\[161\]\[0\] _05863_ _05864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_258_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_157_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15278_ _00036_ net4 mod.u_scanchain_local.module_data_in\[35\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_89_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_208_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14229_ _00083_ net3 mod.u_cpu.rf_ram.memory\[573\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_176_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11535__A1 _05164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_193_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12583__I0 _05869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08400__A1 _01709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_217_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10091__I _04136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_258_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09770_ _03936_ mod.u_cpu.rf_ram.memory\[551\]\[1\] _03943_ _03947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_101_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13288__A1 _06377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14734__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_67_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08721_ _02591_ _03020_ _03027_ _01657_ _03028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__13827__A3 _06643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11915__I _05405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08703__A2 _02999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13108__S _06239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09900__A1 _03837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08652_ _02136_ _02958_ _02959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_39_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_82_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07603_ _01891_ _01901_ _01910_ _01911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_54_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08583_ _01722_ mod.u_cpu.rf_ram.memory\[286\]\[1\] _02889_ _02030_ _02890_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__14884__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07534_ mod.u_cpu.rf_ram.memory\[320\]\[0\] mod.u_cpu.rf_ram.memory\[321\]\[0\] mod.u_cpu.rf_ram.memory\[322\]\[0\]
+ mod.u_cpu.rf_ram.memory\[323\]\[0\] _01841_ _01763_ _01842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_179_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_223_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08467__A1 _02303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_223_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_224_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07465_ _01750_ _01773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_210_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09204_ mod.u_arbiter.i_wb_cpu_rdt\[27\] mod.u_arbiter.i_wb_cpu_dbus_dat\[24\] _03474_
+ _03475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_139_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07396_ _01538_ _01704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_241_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11074__I0 _04841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09135_ mod.u_arbiter.i_wb_cpu_dbus_dat\[0\] _03430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_202_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10266__I _04248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09066_ _03361_ _03368_ _03369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_194_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14264__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08017_ _02109_ _02325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_150_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13515__A2 _06568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_265_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07508__C _01815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09968_ _03919_ _04087_ _04088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_89_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08919_ mod.u_cpu.rf_ram.memory\[536\]\[1\] mod.u_cpu.rf_ram.memory\[537\]\[1\] mod.u_cpu.rf_ram.memory\[538\]\[1\]
+ mod.u_cpu.rf_ram.memory\[539\]\[1\] _02560_ _02495_ _03226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_4225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_170_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09899_ _04041_ _00161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_92_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11930_ _05436_ _00797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_58_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_217_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_206_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11861_ _05386_ _05387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13600_ _03713_ _04922_ _06621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_2856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10812_ _04668_ _04669_ _04670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_260_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08458__A1 _02759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14580_ _00434_ net3 mod.u_cpu.rf_ram.memory\[397\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11792_ mod.u_cpu.rf_ram.memory\[233\]\[0\] _04954_ _05339_ _05340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_129_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_213_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13531_ _06582_ _01252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_10743_ _04574_ _04623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_201_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_201_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_13462_ _03569_ _06531_ _06532_ _03574_ _06535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_201_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13203__A1 _06118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10674_ _04577_ _00400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_199_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_15201_ _01054_ net3 mod.u_cpu.rf_ram.memory\[137\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_127_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12413_ _05761_ mod.u_cpu.rf_ram.memory\[175\]\[1\] _05758_ _05762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_103_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__14607__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_185_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13393_ _06442_ _06398_ _06486_ _06487_ _06488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__11765__A1 _04377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15132_ _00985_ net3 mod.u_cpu.rf_ram.memory\[166\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12344_ _05715_ _00932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08630__A1 _02097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15063_ _00917_ net3 mod.u_cpu.rf_ram.memory\[188\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__13506__A2 _03250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10904__I _03803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12275_ _04984_ _05668_ _05669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11517__A1 _04732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14757__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_175_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14014_ mod.u_arbiter.i_wb_cpu_dbus_dat\[17\] _06966_ _06973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11226_ _04952_ mod.u_cpu.rf_ram.memory\[326\]\[1\] _04949_ _04953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_136_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_218_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11936__S _05439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11157_ _04360_ _04906_ _04907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_67_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10108_ _04043_ _04186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_95_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11088_ _04859_ _04848_ _04860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_5471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_114_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_264_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10879__I0 _04698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14916_ _00770_ net3 mod.u_cpu.rf_ram.memory\[228\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10039_ _04136_ _04137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_82_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08697__A1 _02204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13690__A1 _06693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08249__C _02491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14847_ _00701_ net3 mod.u_cpu.rf_ram.memory\[264\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_84_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_263_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_252_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_205_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08449__A1 _02337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_14778_ _00632_ net3 mod.u_cpu.rf_ram.memory\[298\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_264_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08839__I3 _03145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_205_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13729_ _06429_ _06732_ _06734_ _06735_ _06736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_232_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11470__I _05119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_176_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07250_ _01511_ _01557_ _01558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_32_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13045__I1 mod.u_cpu.rf_ram.memory\[107\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_223_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14287__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11056__I0 _04825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15532__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07181_ _01488_ _01489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_185_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09875__I _04024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_219_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07395__I _01702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_160_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13902__C1 _06699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09822_ _03985_ _03986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_63_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_259_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_228_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09753_ _03932_ _03933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_230_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08704_ _01486_ _03010_ _03011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__14021__I _06942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08688__A1 _02179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09684_ _03809_ _03878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_254_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_215_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09115__I _03413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08635_ _02097_ _02941_ _02942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_265_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12677__S _05941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07360__A1 _01662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_242_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15062__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08566_ _01791_ _02863_ _02872_ _02873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_223_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07517_ _01743_ _01825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_120_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08535__S1 _01916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08497_ _02672_ _02803_ _02804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_211_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07448_ _01728_ mod.u_cpu.rf_ram.memory\[420\]\[0\] _01755_ _01756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_211_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07663__A2 mod.u_cpu.rf_ram.memory\[302\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08860__A1 _01468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07379_ _01686_ _01687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_148_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_202_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09118_ _03413_ _03417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_129_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10390_ _04365_ mod.u_cpu.rf_ram.memory\[460\]\[0\] _04385_ _04386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_109_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_191_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_198_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09049_ _03352_ mod.u_cpu.cpu.o_wdata0 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_191_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12060_ _05523_ _00840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_172_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12172__A1 _05325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11011_ _04806_ _00508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_137_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4000 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4011 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_77_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4022 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4033 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_213_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4044 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4055 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12962_ _06138_ _06139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4066 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15405__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4077 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_218_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4088 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11913_ _05413_ mod.u_cpu.rf_ram.memory\[223\]\[0\] _05424_ _05425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_3343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14701_ _00555_ net3 mod.u_cpu.rf_ram.memory\[337\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_4099 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_248_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_245_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12893_ _06073_ mod.u_cpu.rf_ram.memory\[98\]\[0\] _06084_ _06085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_234_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11844_ _05366_ mod.u_cpu.rf_ram.memory\[159\]\[0\] _05375_ _05376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_14632_ _00486_ net3 mod.u_cpu.rf_ram.memory\[371\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_261_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1930 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1941 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_202_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1952 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_14563_ _00417_ net3 mod.u_cpu.rf_ram.memory\[406\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1963 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11775_ _05106_ _05328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__15555__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11290__I _04951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1974 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_158_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1985 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1996 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10726_ _04611_ _04610_ _04612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_13514_ mod.u_cpu.cpu.state.o_cnt_r\[1\] _03388_ _03337_ _06568_ _06569_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_14494_ _00348_ net3 mod.u_cpu.rf_ram.memory\[440\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_13445_ _06524_ _01224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_173_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10657_ _04290_ _04437_ _04565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_220_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11738__A1 _05300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11589__I1 mod.u_cpu.rf_ram.memory\[268\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12786__I0 _05998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13376_ _06130_ _06472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_126_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10588_ _04518_ _00373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_103_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15115_ _00968_ net3 mod.u_cpu.rf_ram.memory\[419\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12327_ _05667_ _05703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_103_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15046_ _00900_ net3 mod.u_cpu.rf_ram.memory\[196\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12258_ _05656_ _00905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_141_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_218_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11209_ _04941_ _00571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_253_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12189_ _05609_ mod.u_cpu.rf_ram.memory\[203\]\[1\] _05607_ _05610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_190_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10713__A2 _04570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_231_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15085__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_114_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13663__A1 _06661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtiny_user_project_160 wbs_dat_o[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_97_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12466__A2 _05803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_236_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__12710__I0 _05963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtiny_user_project_171 wbs_dat_o[21] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_209_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07342__A1 _01643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08420_ mod.u_cpu.rf_ram.memory\[415\]\[1\] _02727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_224_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07893__A2 _02199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_229_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10229__A1 _04272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_251_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08351_ _02085_ mod.u_cpu.rf_ram.memory\[492\]\[1\] _02658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_260_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07302_ _01608_ _01609_ _01610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_149_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08282_ _02560_ _02587_ _02588_ _02188_ _02589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_220_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14215__I0 _03735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14922__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_177_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08842__A1 _02272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_220_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07233_ mod.u_cpu.rf_ram.memory\[456\]\[0\] mod.u_cpu.rf_ram.memory\[457\]\[0\] mod.u_cpu.rf_ram.memory\[458\]\[0\]
+ mod.u_cpu.rf_ram.memory\[459\]\[0\] _01540_ _01501_ _01541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__13718__A2 _06123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_192_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12777__I0 _05992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07164_ _01462_ mod.u_cpu.cpu.immdec.imm19_12_20\[6\] _01473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_117_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10401__A1 _04242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08070__A2 _02368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12529__I0 _05837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14302__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07853__I _01646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15428__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09805_ _03856_ _03966_ _03973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_75_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07997_ _02303_ _02304_ _02305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_87_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07581__A1 _01849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_216_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09736_ _03902_ _03919_ _03920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_55_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_255_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_228_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09322__A2 _03538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10468__A1 _03991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09667_ _03864_ _03865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__14452__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_227_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15578__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_216_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07333__A1 _01608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08618_ _01849_ _02924_ _02925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_42_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_243_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09598_ _03802_ mod.u_cpu.rf_ram.memory\[56\]\[0\] _03811_ _03812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12209__A2 _04125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13406__A1 _04223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08549_ mod.u_cpu.rf_ram.memory\[317\]\[1\] _02856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11968__A1 _04025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11560_ _05180_ mod.u_cpu.rf_ram.memory\[273\]\[0\] _05181_ _05182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_51_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_243_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08833__A1 _01592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_196_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10511_ _04467_ mod.u_cpu.rf_ram.memory\[441\]\[1\] _04465_ _04468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_210_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10491__I1 mod.u_cpu.rf_ram.memory\[444\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10640__A1 _04527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11491_ _05135_ _00659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_149_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12768__I0 _05998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_196_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_155_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13230_ _06137_ _06133_ _06337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_10442_ _04277_ _04407_ _04420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_171_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08352__C _02067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_200_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__11440__I0 _05087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_170_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13161_ mod.u_arbiter.i_wb_cpu_rdt\[31\] mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat\[15\]
+ _06268_ _06272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_48_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10373_ _04308_ _04373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_164_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12112_ _05557_ _00858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_156_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13092_ _06204_ _06230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_46_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_85_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12043_ _05511_ _00835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_78_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07247__S1 _01501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07763__I _01746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_250_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11285__I _04988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__12448__A2 _05784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13994_ _06910_ _06958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_93_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_218_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_206_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12945_ _03498_ _06122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_3151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_234_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08808__B _03114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_248_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07875__A2 mod.u_cpu.rf_ram.memory\[206\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12876_ _05494_ _05263_ _06074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__14945__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_233_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_215_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14615_ _00469_ net3 mod.u_cpu.rf_ram.memory\[380\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11827_ _05348_ _05362_ _05363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_2494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15595_ _01366_ net3 mod.u_cpu.rf_ram.memory\[113\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_261_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14070__B2 _07012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_183_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_230_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_159_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11758_ _05187_ _05279_ _05316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_42_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14546_ _00400_ net3 mod.u_cpu.rf_ram.memory\[414\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_92_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_202_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10709_ _04598_ mod.u_cpu.rf_ram.memory\[408\]\[0\] _04600_ _04601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10631__A1 _04414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11689_ _05139_ _05255_ _05269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_186_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14477_ _00331_ net3 mod.u_cpu.rf_ram.memory\[44\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_146_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13428_ _03371_ _06511_ _06514_ _03492_ _06515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_155_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13420__I1 mod.u_cpu.rf_ram.memory\[339\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08262__C _02539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_259_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13359_ _06454_ _06455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_155_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08052__A2 mod.u_cpu.rf_ram.memory\[70\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14325__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_114_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_216_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07920_ _02225_ _02226_ _02227_ _01683_ _02228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_64_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_69_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15029_ _00883_ net3 mod.u_cpu.rf_ram.memory\[203\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_190_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12687__A2 _05947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07673__I _01750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12931__I0 _06105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07851_ _02157_ _02158_ _02159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_25_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14475__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_229_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07563__A1 _01852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xinput2 io_in[11] net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07782_ _01661_ _02090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_256_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_237_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09521_ _03744_ _03745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_209_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07315__A1 _01573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_227_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09452_ mod.u_cpu.cpu.decode.opcode\[1\] _03679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_225_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_225_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_213_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_213_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08403_ _02687_ _02702_ _02709_ _02606_ _02710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_196_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09383_ mod.u_arbiter.i_wb_cpu_dbus_adr\[24\] _03615_ _03621_ _03622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__10870__A1 _04299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08334_ _02638_ mod.u_cpu.rf_ram.memory\[502\]\[1\] _02640_ _01615_ _02641_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_221_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15100__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08265_ mod.u_cpu.rf_ram.memory\[541\]\[0\] _02573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_165_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07216_ _01523_ _01524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08196_ _02455_ _02499_ _02503_ _02467_ _02504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_146_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07147_ mod.u_cpu.cpu.immdec.imm24_20\[1\] _01451_ _01455_ _01456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_106_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15250__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14818__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08426__S0 _02688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_114_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__14968__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09504__S _03729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09719_ _03877_ mod.u_cpu.rf_ram.memory\[556\]\[0\] _03906_ _03907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_216_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10991_ _04791_ _00503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_216_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11833__I _03959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_216_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12730_ _05977_ _01056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_231_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07857__A2 mod.u_cpu.rf_ram.memory\[198\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_204_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09303__I _03495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_215_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_150_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12661_ _05918_ mod.u_cpu.rf_ram.memory\[144\]\[0\] _05931_ _05932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_43_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_248_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_203_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11612_ _05199_ mod.u_cpu.rf_ram.memory\[264\]\[0\] _05215_ _05216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14400_ _00254_ net3 mod.u_cpu.rf_ram.memory\[487\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_70_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_212_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15380_ _01155_ net3 mod.u_cpu.rf_ram.memory\[69\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08806__A1 _02665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12592_ _05885_ _01010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12602__A2 _05882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_156_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_211_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11543_ _05162_ mod.u_cpu.rf_ram.memory\[276\]\[1\] _05168_ _05170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_204_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14331_ _00185_ net3 mod.u_cpu.rf_ram.memory\[522\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_141_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14348__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_184_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07758__I _01704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14262_ _00116_ net3 mod.u_cpu.rf_ram.memory\[556\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11474_ _05108_ mod.u_cpu.rf_ram.memory\[287\]\[1\] _05121_ _05123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09606__I0 _03800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_104_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13213_ _06118_ _06320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_137_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10425_ _04400_ mod.u_cpu.rf_ram.memory\[454\]\[0\] _04408_ _04409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_124_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14193_ _07092_ _05803_ _07093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_152_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13144_ _06262_ _01185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_139_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10356_ _04348_ mod.u_cpu.rf_ram.memory\[465\]\[0\] _04361_ _04362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_152_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14498__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07793__A1 _01836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13075_ _03713_ _05640_ _06219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_254_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10287_ _03781_ _04315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__13866__A1 _06791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12913__I0 _06086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12026_ _05483_ _05501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_266_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07426__C _01529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_211_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_238_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_219_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13977_ _06944_ _06945_ _01335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_93_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12928_ _05742_ _04704_ _06108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_262_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_221_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10852__A1 _04290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15123__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12859_ mod.u_cpu.rf_ram_if.rtrig1 mod.u_cpu.rf_ram.rdata\[1\] _06061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_178_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15578_ _01349_ net3 mod.u_arbiter.i_wb_cpu_dbus_dat\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09845__I0 _04001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_203_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_202_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12574__I _05873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14529_ _00383_ net3 mod.u_cpu.rf_ram.memory\[423\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_187_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_186_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_147_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08273__A2 _02572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08050_ _01823_ _02357_ _02358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__15273__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_190_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11404__I0 _05071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11918__I _03750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13157__I0 mod.u_arbiter.i_wb_cpu_rdt\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08720__C _02347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08952_ _03256_ _03257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_115_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13857__A1 _06487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07903_ _01924_ _02211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__09525__A2 _03747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08883_ _02456_ mod.u_cpu.rf_ram.memory\[572\]\[1\] _03189_ _03190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_57_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07834_ _02110_ _02133_ _02140_ _02141_ _02142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_29_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_217_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3909 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07765_ _02053_ _02072_ _02073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__11653__I _05221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_186_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12132__I1 mod.u_cpu.rf_ram.memory\[208\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09504_ mod.u_cpu.rf_ram.memory\[9\]\[0\] _03699_ _03729_ _03730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_266_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_213_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07696_ _01722_ mod.u_cpu.rf_ram.memory\[286\]\[0\] _02003_ _01970_ _02004_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__10143__I0 _04193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_164_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09435_ mod.u_cpu.cpu.immdec.imm11_7\[0\] mod.u_cpu.cpu.immdec.imm11_7\[1\] _03664_
+ _03665_ _03666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_73_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_252_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_197_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14034__A1 mod.u_arbiter.i_wb_cpu_rdt\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_36_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09366_ _03605_ _03606_ _03607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__15616__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_240_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12596__A1 _05888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08317_ mod.u_cpu.rf_ram.memory\[471\]\[1\] _02624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_21_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11643__I0 _05222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09461__A1 _03681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09297_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[11\] mod.u_cpu.cpu.ctrl.o_ibus_adr\[10\] _03543_
+ _03549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_227_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_201_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08248_ _02545_ _02549_ _02554_ _02555_ _02556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_123_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10071__A2 _04143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_197_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_197_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14640__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_181_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08179_ _02010_ _02487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_107_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08647__S0 _02125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09793__I _03889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12899__A2 _06048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10210_ _04186_ _04259_ _04260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_180_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11190_ _04916_ mod.u_cpu.rf_ram.memory\[332\]\[1\] _04927_ _04929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08567__A3 _02873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11571__A2 _05188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13148__I0 mod.u_arbiter.i_wb_cpu_rdt\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10141_ _03872_ _04209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_121_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14790__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10072_ _04148_ mod.u_cpu.rf_ram.memory\[506\]\[0\] _04159_ _04160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_251_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_198_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07527__A1 _01818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_102_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12520__A1 _05355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_153_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13900_ _06677_ _06885_ _01318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_48_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_248_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14880_ _00734_ net3 mod.u_cpu.rf_ram.memory\[243\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_208_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_262_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13831_ _06135_ _06826_ _06828_ _01306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_75_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15146__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12123__I1 mod.u_cpu.rf_ram.memory\[20\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_90_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_204_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10974_ _04227_ _04779_ _04780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_13762_ _03298_ mod.u_cpu.cpu.immdec.imm24_20\[0\] _06421_ _06766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__10134__I0 _04199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_250_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_244_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_216_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_15501_ _01272_ net3 mod.u_arbiter.i_wb_cpu_dbus_adr\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_203_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12713_ _05966_ mod.u_cpu.rf_ram.memory\[7\]\[1\] _05964_ _05967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_15_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10834__A1 _04277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_188_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13693_ mod.u_cpu.cpu.immdec.imm19_12_20\[2\] _06658_ _06700_ _06702_ _06703_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_70_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15432_ _01207_ net3 mod.u_cpu.cpu.immdec.imm11_7\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__15296__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_231_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12644_ _05732_ _05920_ _05921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_19_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_197_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08805__C _01669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12575_ _05874_ mod.u_cpu.rf_ram.memory\[15\]\[1\] _05871_ _05875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_15363_ _01138_ net3 mod.u_cpu.rf_ram.memory\[85\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_200_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_196_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_200_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11004__S _04799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14314_ _00168_ net3 mod.u_cpu.rf_ram.memory\[530\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11526_ _05158_ _00671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_117_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15294_ _00054_ net4 mod.u_scanchain_local.module_data_in\[51\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_7_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11457_ _05110_ _03782_ _05111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_14245_ _00099_ net3 mod.u_cpu.rf_ram.memory\[565\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10843__S _04688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08638__S0 _02106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13000__A2 _06166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10408_ mod.u_cpu.rf_ram.memory\[457\]\[0\] _04396_ _04397_ _04398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_139_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14176_ _07082_ _01397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_11388_ _04531_ _05065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_152_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13139__I0 mod.u_arbiter.i_wb_cpu_rdt\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13127_ _06252_ _06253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_10339_ _04350_ _00292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_97_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09507__A2 _03352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13058_ _06208_ _01153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_140_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12009_ _05484_ mod.u_cpu.rf_ram.memory\[575\]\[1\] _05486_ _05490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_266_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_254_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_266_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08810__S0 _02366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08191__A1 _02456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_187_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07550_ _01758_ _01858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_228_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_207_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14513__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15639__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12814__A2 _06031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_146_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_234_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_179_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07481_ _01770_ _01772_ _01786_ _01788_ _01789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_185_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09220_ _03410_ mod.u_scanchain_local.module_data_in\[36\] _03484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07900__B _02207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_210_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_166_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14663__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09151_ mod.u_arbiter.i_wb_cpu_rdt\[6\] _03441_ _03442_ _03443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10428__I1 mod.u_cpu.rf_ram.memory\[454\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_187_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08102_ _01646_ _02410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_124_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11250__A1 _04831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09082_ net1 _03383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_148_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08033_ _01696_ _02340_ _02321_ _02341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_162_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15019__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08629__S0 _02085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07757__A1 _01849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12750__A1 _02162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_130_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09984_ _04091_ mod.u_cpu.rf_ram.memory\[520\]\[1\] _04097_ _04099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_192_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09118__I _03413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08935_ _02545_ _03238_ _03241_ _02555_ _03242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_131_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15169__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07509__A1 _01656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_170_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08866_ _02462_ _03172_ _03173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_3706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_244_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07817_ _01672_ _02125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__12479__I _05694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08797_ _02348_ _03103_ _01618_ _03104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_85_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_260_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09989__S _04100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07748_ _02053_ _02055_ _02056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_232_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11864__I0 _05385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07679_ _01938_ mod.u_cpu.rf_ram.memory\[278\]\[0\] _01986_ _01952_ _01987_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__14007__A1 _03456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__14007__B2 mod.u_arbiter.i_wb_cpu_dbus_dat\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_198_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09788__I _03959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_201_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_213_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09418_ mod.u_arbiter.i_wb_cpu_dbus_adr\[29\] _03615_ _03651_ _03652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_201_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10690_ _04457_ _04575_ _04588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_41_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08625__C _02077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_178_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09349_ _03588_ _03590_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[19\] _03593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__13230__A2 _06133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_201_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_194_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12360_ _05725_ _05726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11092__I1 mod.u_cpu.rf_ram.memory\[348\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_240_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11311_ _05007_ mod.u_cpu.rf_ram.memory\[313\]\[0\] _05012_ _05013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_194_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_14_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12291_ _05604_ _05679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_113_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14030_ mod.u_arbiter.i_wb_cpu_rdt\[20\] _06976_ _06982_ mod.u_arbiter.i_wb_cpu_dbus_dat\[20\]
+ _06985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_11242_ _04964_ _00581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_84_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08096__S1 _02367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08796__I0 mod.u_cpu.rf_ram.memory\[72\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11173_ _04917_ _00559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_49_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10124_ _04193_ mod.u_cpu.rf_ram.memory\[4\]\[0\] _04197_ _04198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_110_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_212_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14932_ _00786_ net3 mod.u_cpu.rf_ram.memory\[226\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10055_ _04013_ _03859_ _04149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_249_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14536__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4930 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_102_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4941 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_180_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08173__A1 _02479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_263_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_209_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4952 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4963 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14863_ _00717_ net3 mod.u_cpu.rf_ram.memory\[257\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_169_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_4974 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13049__A2 _06201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_247_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4985 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_180_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07920__A1 _02225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4996 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13814_ _06810_ _06813_ _01304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_169_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14794_ _00648_ net3 mod.u_cpu.rf_ram.memory\[290\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_251_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07359__S0 _01664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_189_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_216_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__14686__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13745_ _06656_ _06750_ _06751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_90_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10957_ _04768_ _00492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_44_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_56_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09698__I _03762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10283__A2 _04310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13676_ _06437_ _06448_ _06686_ _06372_ _06687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_10888_ _04389_ _04108_ _04722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_148_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13757__B1 _06713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15415_ _01190_ net3 mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_12627_ _05904_ mod.u_cpu.rf_ram.memory\[150\]\[0\] _05909_ _05910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XPHY_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08079__I2 mod.u_cpu.rf_ram.memory\[2\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09425__A1 mod.u_arbiter.i_wb_cpu_dbus_adr\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_157_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10035__A2 _03715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08107__I _01765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15346_ _01121_ net3 mod.u_cpu.rf_ram.memory\[389\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_200_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12558_ _05657_ _05757_ _05863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07531__S0 _01837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11509_ _05147_ mod.u_cpu.rf_ram.memory\[282\]\[1\] _05145_ _05148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_145_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12852__I _03398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15277_ _00035_ net4 mod.u_scanchain_local.module_data_in\[34\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12489_ _05807_ mod.u_cpu.rf_ram.memory\[171\]\[1\] _05817_ _05819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_176_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14228_ _00082_ net3 mod.u_cpu.rf_ram.memory\[573\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12032__I0 _05501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_217_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_259_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11535__A2 _05130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12732__A1 _03932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15311__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_193_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_140_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14159_ _06153_ _03270_ _01407_ _07070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_98_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_256_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_113_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_224_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08720_ _01698_ _03023_ _03026_ _02347_ _03027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__09382__B _03417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_227_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_255_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07681__I _01886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15461__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_226_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08651_ mod.u_cpu.rf_ram.memory\[167\]\[1\] _02958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_67_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09900__A2 _04033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_227_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07911__A1 _01607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_242_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07602_ _01872_ _01902_ _01909_ _01657_ _01910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_82_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08582_ _02027_ _02888_ _02889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_214_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07533_ _01710_ _01841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_241_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__11846__I0 _05364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11931__I _03698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_179_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_179_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11471__A1 _04700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07464_ mod.u_cpu.rf_ram.memory\[424\]\[0\] mod.u_cpu.rf_ram.memory\[425\]\[0\] mod.u_cpu.rf_ram.memory\[426\]\[0\]
+ mod.u_cpu.rf_ram.memory\[427\]\[0\] _01753_ _01771_ _01772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_179_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09203_ _03414_ _03474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_07395_ _01702_ _01703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_72_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_210_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_202_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_194_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09134_ _03428_ _03387_ _03421_ _03429_ _00063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_148_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08017__I _02109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_198_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07978__A1 _02129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14409__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12762__I _05937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09065_ _03300_ _03367_ _03368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07856__I _01820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_190_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08016_ mod.u_cpu.rf_ram.memory\[112\]\[0\] mod.u_cpu.rf_ram.memory\[113\]\[0\] mod.u_cpu.rf_ram.memory\[114\]\[0\]
+ mod.u_cpu.rf_ram.memory\[115\]\[0\] _01664_ _02323_ _02324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_151_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_194_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11378__I _04995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08180__C _02487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_235_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10585__I0 _04506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14559__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_249_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09967_ _03995_ _04087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_4204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_218_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_170_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08918_ _03215_ _03224_ _01447_ _03225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_4226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09898_ _04036_ mod.u_cpu.rf_ram.memory\[534\]\[1\] _04039_ _04041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_4237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_218_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08849_ _03001_ _03155_ _03156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_3525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_206_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_261_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11860_ _03726_ _04378_ _05386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_2824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_214_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11837__I0 _05364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10811_ _04569_ _04669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_11791_ _05078_ _05320_ _05339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_2868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_198_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08458__A2 _02760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11841__I _05372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_198_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13530_ _06581_ mod.u_cpu.rf_ram.memory\[129\]\[1\] _06579_ _06582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_198_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10742_ _04621_ _04622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_41_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_230_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_139_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13461_ _06534_ _01230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__10457__I _04429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10673_ _04557_ mod.u_cpu.rf_ram.memory\[414\]\[0\] _04576_ _04577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__13203__A2 _06309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15200_ _01053_ net3 mod.u_cpu.rf_ram.memory\[137\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_167_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12412_ _05710_ _05761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_138_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13392_ _06470_ _06397_ _06487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_139_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_194_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07969__A1 _01742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_182_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11765__A2 _05320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15131_ _00984_ net3 mod.u_cpu.rf_ram.memory\[167\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__15334__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12343_ _05713_ mod.u_cpu.rf_ram.memory\[182\]\[0\] _05714_ _05715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_181_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08630__A2 _02936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12014__I0 _05484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15062_ _00916_ net3 mod.u_cpu.rf_ram.memory\[188\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12274_ _05667_ _05668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_182_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_253_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11225_ _04951_ _04952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_14013_ _06969_ _06972_ _01344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_4_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__15484__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11156_ _04905_ _04906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08784__I3 mod.u_cpu.rf_ram.memory\[87\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10107_ _04184_ _04173_ _04185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_136_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_191_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11087_ _03780_ _04859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_237_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_208_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14915_ _00769_ net3 mod.u_cpu.rf_ram.memory\[39\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10038_ _04135_ _04136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_76_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08697__A2 mod.u_cpu.rf_ram.memory\[196\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13690__A2 _06463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_224_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_4782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14846_ _00700_ net3 mod.u_cpu.rf_ram.memory\[264\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_4793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_223_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14777_ _00631_ net3 mod.u_cpu.rf_ram.memory\[2\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_16_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08449__A2 _02755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11989_ _02485_ _05475_ _05476_ _00816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_182_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13728_ _06494_ _06735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_108_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_225_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_225_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07752__S0 _02059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_182_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13659_ _06371_ _06670_ _06671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_143_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_220_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11205__A1 _04808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_176_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07180_ _01487_ _01488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_34_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_118_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_258_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_158_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12953__A1 _06125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15329_ mod.u_cpu.cpu.o_wen1 net3 mod.u_cpu.rf_ram_if.wen1_r vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_173_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14701__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13902__B1 _06693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13902__C2 _06135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_232_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_235_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09821_ _03984_ _03985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_99_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14851__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09752_ _03931_ _03932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_100_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08137__A1 _02337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09334__B1 _03555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_227_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08703_ _02997_ _02999_ _01891_ _03009_ _03010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_100_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09683_ _03739_ _03877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07344__C _01651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08688__A2 mod.u_cpu.rf_ram.memory\[204\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_243_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__15207__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08634_ mod.u_cpu.rf_ram.memory\[188\]\[1\] mod.u_cpu.rf_ram.memory\[189\]\[1\] mod.u_cpu.rf_ram.memory\[190\]\[1\]
+ mod.u_cpu.rf_ram.memory\[191\]\[1\] _02092_ _02098_ _02941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_215_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07360__A2 _01667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11819__I0 _05350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08565_ _01956_ _02864_ _02871_ _01989_ _02872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_35_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07516_ mod.u_cpu.rf_ram.memory\[348\]\[0\] mod.u_cpu.rf_ram.memory\[349\]\[0\] mod.u_cpu.rf_ram.memory\[350\]\[0\]
+ mod.u_cpu.rf_ram.memory\[351\]\[0\] _01823_ _01821_ _01824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_08496_ mod.u_cpu.rf_ram.memory\[335\]\[1\] _02803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_126_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12492__I0 _05813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_210_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_195_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14231__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13789__S _03502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07447_ _01753_ _01754_ _01755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__15357__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10277__I _03769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12693__S _05953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_183_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07378_ _01527_ _01686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_129_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12944__A1 _06118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09117_ _03279_ _03416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_164_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14381__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_191_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09048_ _03250_ _03348_ _03351_ _03352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_190_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10558__I0 _04498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11010_ _04803_ mod.u_cpu.rf_ram.memory\[360\]\[0\] _04805_ _04806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_78_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12172__A2 _05576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_131_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10740__I _03737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_219_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4001 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4012 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4023 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4034 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_161_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4045 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08210__I _02291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_180_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_12961_ _06137_ _06138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08518__I3 mod.u_cpu.rf_ram.memory\[339\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4056 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4067 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_248_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_206_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4078 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14700_ _00554_ net3 mod.u_cpu.rf_ram.memory\[337\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_4089 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11912_ _04845_ _05423_ _05424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_3344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12892_ _03974_ _06048_ _06084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_3366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_205_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14631_ _00485_ net3 mod.u_cpu.rf_ram.memory\[372\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_72_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11843_ _04845_ _05374_ _05375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_260_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_221_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1920 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_199_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_214_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1942 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_199_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_214_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_199_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14562_ _00416_ net3 mod.u_cpu.rf_ram.memory\[406\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1953 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11774_ _05327_ _00750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1964 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_214_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1975 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08300__A1 _02083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1986 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_202_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13513_ _05791_ _06568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_207_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_186_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1997 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10725_ _04541_ _04611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_186_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14493_ _00347_ net3 mod.u_cpu.rf_ram.memory\[441\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_201_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_186_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14724__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13444_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[7\] _06519_ _06520_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[8\]
+ _06524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_186_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10656_ _04564_ _00395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_103_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__13498__I _06537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12108__S _05553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13375_ _06470_ _06471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_155_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10587_ _04514_ mod.u_cpu.rf_ram.memory\[428\]\[1\] _04516_ _04518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_6_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15114_ _00967_ net3 mod.u_cpu.rf_ram.memory\[419\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_155_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12326_ _05702_ _00927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_86_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_114_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14874__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_181_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15045_ _00899_ net3 mod.u_cpu.rf_ram.memory\[109\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12257_ _05635_ mod.u_cpu.rf_ram.memory\[194\]\[1\] _05654_ _05656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_5_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08367__A1 _02672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_214_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11208_ _04936_ mod.u_cpu.rf_ram.memory\[32\]\[1\] _04939_ _04941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_12188_ _05549_ _05609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_64_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_123_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_214_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_95_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_256_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11139_ _04883_ mod.u_cpu.rf_ram.memory\[340\]\[0\] _04894_ _04895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_95_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_209_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_49_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xtiny_user_project_150 wbs_dat_o[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_48_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xtiny_user_project_161 wbs_dat_o[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_3_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xtiny_user_project_172 wbs_dat_o[22] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_225_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12710__I1 mod.u_cpu.rf_ram.memory\[7\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_252_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07342__A2 mod.u_cpu.rf_ram.memory\[494\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14254__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14829_ _00683_ net3 mod.u_cpu.rf_ram.memory\[273\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_36_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11481__I _05107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_224_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10229__A2 _04263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08350_ mod.u_cpu.rf_ram.memory\[493\]\[1\] _02657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__11426__A1 _04812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_189_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07301_ mod.u_cpu.rf_ram.memory\[509\]\[0\] _01609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_220_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08281_ _02198_ mod.u_cpu.rf_ram.memory\[460\]\[1\] _02588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08842__A2 mod.u_cpu.rf_ram.memory\[44\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13179__A1 _06122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_177_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07232_ _01539_ _01540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_160_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07163_ mod.u_cpu.cpu.immdec.imm24_20\[2\] _01467_ _01472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_9_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_191_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_236_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_259_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09804_ _03972_ _00135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_86_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07996_ mod.u_cpu.rf_ram.memory\[111\]\[0\] _02304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_75_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09735_ _03918_ _03919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_74_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_228_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10468__A2 _04437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09666_ _03768_ _03848_ _03864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_216_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_35 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08617_ mod.u_cpu.rf_ram.memory\[136\]\[1\] mod.u_cpu.rf_ram.memory\[137\]\[1\] mod.u_cpu.rf_ram.memory\[138\]\[1\]
+ mod.u_cpu.rf_ram.memory\[139\]\[1\] _02022_ _02043_ _02924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_242_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09597_ _03805_ _03810_ _03811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08548_ mod.u_cpu.rf_ram.memory\[312\]\[1\] mod.u_cpu.rf_ram.memory\[313\]\[1\] mod.u_cpu.rf_ram.memory\[314\]\[1\]
+ mod.u_cpu.rf_ram.memory\[315\]\[1\] _01802_ _01932_ _02855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__14747__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_208_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_211_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08479_ _01997_ _02782_ _02785_ _02096_ _02786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__12217__I0 _05609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10510_ _04429_ _04467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_11490_ _05128_ mod.u_cpu.rf_ram.memory\[285\]\[1\] _05131_ _05135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_13_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10640__A2 _04389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14897__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10441_ _04419_ _00325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_109_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08597__A1 _02070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13160_ _06271_ _01192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_10372_ _04372_ _00303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11440__I1 mod.u_cpu.rf_ram.memory\[292\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_191_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_191_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12111_ _05539_ mod.u_cpu.rf_ram.memory\[68\]\[0\] _05556_ _05557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_163_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13091_ _06229_ _01165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_152_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_105_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12042_ _05501_ mod.u_cpu.rf_ram.memory\[60\]\[1\] _05509_ _05511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__13342__A1 _06438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_254_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_266_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12940__I1 mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_266_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_238_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_266_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_219_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14142__I0 _07055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_266_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14277__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_265_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_13993_ mod.u_arbiter.i_wb_cpu_dbus_dat\[12\] _06954_ _06957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09849__A1 _03771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15522__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_207_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12944_ _06118_ _06120_ _06121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_3141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08521__A1 _01893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08808__C _02380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_206_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_222_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12875_ _06072_ _06073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_261_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_209_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_234_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14614_ _00468_ net3 mod.u_cpu.rf_ram.memory\[380\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11826_ _04294_ _03942_ _05362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15594_ _01365_ net3 mod.u_cpu.rf_ram.memory\[113\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14545_ _00399_ net3 mod.u_cpu.rf_ram.memory\[415\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11757_ _05315_ _00745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_187_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10708_ _04168_ _04599_ _04600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10631__A2 _04548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14476_ _00330_ net3 mod.u_cpu.rf_ram.memory\[44\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11688_ _05221_ _05268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_179_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_220_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08543__C _01504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10645__I _04522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13427_ _06513_ _06514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_179_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_139_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10639_ _04553_ _00389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_127_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13358_ _06395_ _06380_ _06131_ _06454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_154_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10395__A1 _03727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_255_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_170_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12309_ _05679_ mod.u_cpu.rf_ram.memory\[185\]\[0\] _05690_ _05691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_115_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15052__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13289_ _03501_ _03428_ _06386_ _06387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_142_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13333__A1 _06318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09147__S _03439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15028_ _00882_ net3 mod.u_cpu.rf_ram.memory\[203\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_130_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10147__A1 _04068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11476__I _05118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_190_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13884__A2 _06311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07850_ mod.u_cpu.rf_ram.memory\[197\]\[0\] _02158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_257_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_190_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08760__A1 _02631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07563__A2 _01853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14133__I0 _07043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_232_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07781_ _01818_ _02082_ _02088_ _02089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
Xinput3 io_in[12] net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_20
XFILLER_110_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09520_ _03741_ _03743_ _03744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_49_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_225_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_213_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09451_ _03678_ _03294_ _03677_ _00006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_224_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_197_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08402_ _02654_ _02705_ _02708_ _01979_ _02709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_09382_ _03564_ _03617_ _03620_ _03417_ _03621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XANTENNA__10870__A2 _04709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_240_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08333_ _02197_ _02639_ _02640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_127_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_220_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08264_ mod.u_cpu.rf_ram.memory\[536\]\[0\] mod.u_cpu.rf_ram.memory\[537\]\[0\] mod.u_cpu.rf_ram.memory\[538\]\[0\]
+ mod.u_cpu.rf_ram.memory\[539\]\[0\] _02450_ _02451_ _02572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_123_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_165_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_137_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07215_ _01497_ _01523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10555__I _03761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08195_ _02461_ mod.u_cpu.rf_ram.memory\[574\]\[0\] _02502_ _02465_ _02503_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_203_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_193_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08579__A1 _01711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_119_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07146_ _01452_ _01454_ _01448_ _01425_ _01455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_69_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_192_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_173_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_238_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07864__I _01614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08426__S1 _02475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15545__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08751__A1 _01670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_247_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07979_ mod.u_cpu.rf_ram.memory\[103\]\[0\] _02287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_142_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_216_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_210_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09718_ _03902_ _03905_ _03906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_132_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07813__B _02119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10990_ _04772_ mod.u_cpu.rf_ram.memory\[363\]\[1\] _04789_ _04791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08503__A1 _01520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_216_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09649_ _03850_ _03851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_76_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_243_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_203_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12660_ _05300_ _05920_ _05931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_70_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12438__I0 _05753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_93_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11611_ _04804_ _05214_ _05215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_169_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12063__A1 _04983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12945__I _03498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_208_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_169_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08806__A2 _03105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12591_ _05874_ mod.u_cpu.rf_ram.memory\[156\]\[1\] _05883_ _05885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_243_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_211_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14330_ _00184_ net3 mod.u_cpu.rf_ram.memory\[522\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11542_ _05169_ _00676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_196_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11810__A1 _04808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_221_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_167_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14261_ _00115_ net3 mod.u_cpu.rf_ram.memory\[557\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07490__A1 _01689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11473_ _02002_ _05121_ _05122_ _00654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__15075__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08114__S0 _02421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13212_ _06318_ _06319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_136_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10424_ _04262_ _04407_ _04408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_152_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14192_ mod.u_cpu.rf_ram_if.rgnt _07092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_100_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13143_ mod.u_arbiter.i_wb_cpu_rdt\[23\] mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat\[7\]
+ _06258_ _06262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_10355_ _04360_ _04353_ _04361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_87_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_124_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10286_ _04314_ _00275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13074_ _06218_ _01159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_112_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_219_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13866__A2 _06672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_250_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12025_ _05500_ _00828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11877__A1 _05348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_239_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14912__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08742__A1 _01848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_266_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_266_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_226_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_207_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_266_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11629__A1 _05226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_150_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12677__I0 _05938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13976_ mod.u_arbiter.i_wb_cpu_rdt\[6\] _06938_ _06928_ mod.u_arbiter.i_wb_cpu_dbus_dat\[6\]
+ _06945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_59_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09542__I0 _03764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_202_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12927_ _06072_ _06107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_206_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_111_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_234_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15646_ _01417_ net3 mod.u_cpu.rf_ram.memory\[249\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_222_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12858_ mod.u_cpu.rf_ram_if.rdata1 _06060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_2270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10852__A2 _04687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_181_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_178_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_261_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_203_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11809_ _05351_ _00761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_178_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15577_ _01348_ net3 mod.u_arbiter.i_wb_cpu_dbus_dat\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12789_ _06010_ mod.u_cpu.rf_ram.memory\[130\]\[0\] _06015_ _06016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_221_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_187_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_202_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_230_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15418__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14528_ _00382_ net3 mod.u_cpu.rf_ram.memory\[423\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_147_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_175_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08273__C _02491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13929__I0 _06904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_175_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14459_ _00313_ net3 mod.u_cpu.rf_ram.memory\[458\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_190_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_259_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10368__A1 _04369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14442__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15568__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_192_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_153_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08981__A1 _01428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08951_ _03252_ _03253_ _03255_ _03256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_170_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13857__A2 _06850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07902_ mod.u_cpu.rf_ram.memory\[211\]\[0\] _02210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__11868__A1 _05343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08882_ _02457_ _03188_ _03189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__14592__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_233_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_243_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_229_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07833_ _01716_ _02141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_97_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15553__D _01324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_256_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07764_ mod.u_cpu.rf_ram.memory\[140\]\[0\] mod.u_cpu.rf_ram.memory\[141\]\[0\] mod.u_cpu.rf_ram.memory\[142\]\[0\]
+ mod.u_cpu.rf_ram.memory\[143\]\[0\] _02070_ _02071_ _02072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_09503_ _03714_ _03728_ _03729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_53_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07695_ _01967_ _02002_ _02003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11340__I0 _05032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08592__S0 _01802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_198_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09434_ mod.u_cpu.cpu.immdec.imm11_7\[4\] _03665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_25_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_53_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14034__A2 _06987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_213_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__12045__A1 _05488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09365_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[21\] mod.u_cpu.cpu.ctrl.o_ibus_adr\[20\] _03595_
+ _03606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_178_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15098__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_221_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13793__A1 _06779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08316_ _02566_ mod.u_cpu.rf_ram.memory\[468\]\[1\] _02622_ _02623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__12596__A2 _05882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_240_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09296_ _03541_ _03543_ _03548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__12840__I0 _06035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_177_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09461__A2 _03679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08247_ _02308_ _02555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_119_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_203_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08178_ _02484_ _02485_ _02486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_137_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08647__S1 _02127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07129_ _01425_ _01432_ _01437_ _01438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_238_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08811__I2 mod.u_cpu.rf_ram.memory\[2\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14935__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10140_ _04208_ _00235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08972__A1 _03268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13848__A2 mod.u_arbiter.i_wb_cpu_rdt\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12005__I _03773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10071_ _03797_ _04143_ _04159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_43_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_251_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07527__A2 _01834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12520__A2 _05831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10531__A1 _01793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13830_ mod.u_cpu.cpu.immdec.imm30_25\[4\] _06773_ _06812_ mod.u_cpu.cpu.immdec.imm30_25\[5\]
+ _06827_ _06339_ _06828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_229_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_210_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_260_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_13761_ _03686_ _06764_ _06765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_216_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10973_ _03663_ _04223_ _03724_ _04779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_56_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_262_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_249_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11780__S _05331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15500_ _01271_ net3 mod.u_arbiter.i_wb_cpu_dbus_adr\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__14315__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12712_ _05937_ _05966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__10834__A2 _04669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_204_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13692_ _06656_ _06701_ _06702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_188_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_231_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_204_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15431_ _01206_ net3 mod.u_cpu.cpu.immdec.imm11_7\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_102_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12643_ _05919_ _05920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_31_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_203_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07769__I _01677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_231_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13784__A1 _06065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_15362_ _01137_ net3 mod.u_cpu.rf_ram.memory\[86\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_180_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11634__I1 _05230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12831__I0 _06035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12574_ _05873_ _05874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_156_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08093__C _02361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__14465__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14313_ _00167_ net3 mod.u_cpu.rf_ram.memory\[531\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11525_ _05147_ mod.u_cpu.rf_ram.memory\[27\]\[1\] _05156_ _05158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_156_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10195__I _04248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15293_ _00053_ net4 mod.u_scanchain_local.module_data_in\[50\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_172_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_200_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14244_ _00098_ net3 mod.u_cpu.rf_ram.memory\[565\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_8_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11456_ _04195_ _05110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_172_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08638__S1 _02127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08821__C _01830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10407_ _03714_ _04380_ _04397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_256_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_14175_ _07081_ mod.u_cpu.rf_ram.memory\[88\]\[1\] _07079_ _07082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_217_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11387_ _01964_ _05063_ _05064_ _00626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_98_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13139__I1 mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_180_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13126_ _05785_ _06252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_112_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10338_ _04348_ mod.u_cpu.rf_ram.memory\[468\]\[0\] _04349_ _04350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13839__A2 _06834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13057_ _06199_ mod.u_cpu.rf_ram.memory\[82\]\[1\] _06206_ _06208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_191_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10269_ _04132_ _04300_ _04301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_117_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08715__A1 _02027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12008_ _02501_ _05486_ _05489_ _00822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_121_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08810__S1 _02383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_266_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_238_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08191__A2 mod.u_cpu.rf_ram.memory\[572\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_254_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_207_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12275__A1 _04984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_207_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13959_ _06920_ _05794_ _06930_ _06931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__12786__S _06012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13472__B1 _06540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_207_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_207_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07480_ _01787_ _01788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__15240__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_62_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14808__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15629_ _01400_ net3 mod.u_cpu.rf_ram.memory\[279\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_250_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09818__I1 _03929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_203_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09150_ _03417_ _03442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__10589__A1 _04238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_187_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08101_ _02316_ mod.u_cpu.rf_ram.memory\[20\]\[0\] _02408_ _02409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_159_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15390__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11250__A2 _04969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09081_ _03301_ _03378_ _03382_ _00003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_175_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09894__I _04002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_190_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14958__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08032_ mod.u_cpu.rf_ram.memory\[84\]\[0\] mod.u_cpu.rf_ram.memory\[85\]\[0\] mod.u_cpu.rf_ram.memory\[86\]\[0\]
+ mod.u_cpu.rf_ram.memory\[87\]\[0\] _01857_ _02054_ _02340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_107_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08629__S1 _02086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08731__C _02852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_174_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07206__A1 _01508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10061__I0 _04148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12750__A2 _05989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_192_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09983_ _04098_ _00188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_143_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_192_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08934_ _02550_ mod.u_cpu.rf_ram.memory\[534\]\[1\] _03240_ _02515_ _03241_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_192_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_258_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08865_ mod.u_cpu.rf_ram.memory\[551\]\[1\] _03172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_29_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_218_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07816_ _01687_ _02124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__14338__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_257_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08796_ mod.u_cpu.rf_ram.memory\[72\]\[1\] mod.u_cpu.rf_ram.memory\[73\]\[1\] mod.u_cpu.rf_ram.memory\[74\]\[1\]
+ mod.u_cpu.rf_ram.memory\[75\]\[1\] _02211_ _02386_ _03103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_85_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_226_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07747_ mod.u_cpu.rf_ram.memory\[132\]\[0\] mod.u_cpu.rf_ram.memory\[133\]\[0\] mod.u_cpu.rf_ram.memory\[134\]\[0\]
+ mod.u_cpu.rf_ram.memory\[135\]\[0\] _01893_ _02054_ _02055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_244_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09131__A1 _03424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11864__I1 mod.u_cpu.rf_ram.memory\[70\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07678_ _01949_ _01985_ _01986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_164_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_197_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14007__A2 _06964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14488__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09417_ _03614_ _03649_ _03650_ _03651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_213_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07693__A1 _01998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_244_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11105__S _04870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_240_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_199_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09348_ _03568_ _03591_ _03592_ _00059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_179_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_194_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09279_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[8\] _03533_ _03534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_148_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11310_ _04873_ _05011_ _05012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_154_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_138_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12290_ _05678_ _00915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_165_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11241_ _04952_ mod.u_cpu.rf_ram.memory\[324\]\[1\] _04962_ _04964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10743__I _04574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_1242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_122_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_164_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11172_ _04916_ mod.u_cpu.rf_ram.memory\[335\]\[1\] _04914_ _04917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07257__C _01529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15113__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10123_ _04196_ _03961_ _04197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_5610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14931_ _00785_ net3 mod.u_cpu.rf_ram.memory\[227\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10054_ _04147_ _04148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_94_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_248_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_209_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_4920 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11552__I0 _05159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4931 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_87_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4942 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4953 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14862_ _00716_ net3 mod.u_cpu.rf_ram.memory\[257\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_4964 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15263__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_236_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4975 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_169_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4986 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07920__A2 _02226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13813_ mod.u_cpu.cpu.immdec.imm30_25\[2\] _06773_ _06807_ _06811_ _06812_ mod.u_cpu.cpu.immdec.imm30_25\[3\]
+ _06813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_17_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4997 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14793_ _00647_ net3 mod.u_cpu.rf_ram.memory\[291\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_44_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_250_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_204_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_169_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09122__A1 _03363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_263_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07359__S1 _01666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13744_ mod.u_cpu.cpu.immdec.imm19_12_20\[7\] _06139_ _06338_ _06741_ _06750_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_44_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10956_ _04753_ mod.u_cpu.rf_ram.memory\[368\]\[0\] _04767_ _04768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_147_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13057__I0 _06199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13675_ _06431_ _06490_ _06686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_189_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10887_ _04721_ _00469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_15414_ _01189_ net3 mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_19_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__13757__B2 _06744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12626_ _05494_ _05900_ _05909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_157_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12804__I0 _06019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_197_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09425__A2 _03561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08079__I3 mod.u_cpu.rf_ram.memory\[3\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_200_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15345_ _01120_ net3 mod.u_cpu.rf_ram.memory\[389\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10035__A3 _03717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12557_ _05862_ _00998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_156_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10291__I0 _04313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13509__A1 _06562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11508_ _05107_ _05147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_185_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07531__S1 _01838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15276_ _00034_ net4 mod.u_arbiter.i_wb_cpu_rdt\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12980__A2 _03343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12488_ _05818_ _00973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_144_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11749__I _03696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14182__A1 _03822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14227_ _00081_ net3 mod.u_cpu.rf_ram.memory\[574\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11439_ _05098_ _00644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_172_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08936__A1 _02542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09984__I0 _04091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_14158_ _07069_ _01407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_63_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_152_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13109_ _06241_ _01171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_101_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14089_ _03774_ _07026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_113_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15606__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11543__I0 _05162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11484__I _05119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_239_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08650_ _02129_ mod.u_cpu.rf_ram.memory\[164\]\[1\] _02956_ _02957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_94_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_266_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_266_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_187_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07601_ _01874_ _01905_ _01908_ _01884_ _01909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_255_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08581_ mod.u_cpu.rf_ram.memory\[287\]\[1\] _02888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_82_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_240_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14630__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_226_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_187_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07532_ mod.u_cpu.rf_ram.memory\[340\]\[0\] mod.u_cpu.rf_ram.memory\[341\]\[0\] mod.u_cpu.rf_ram.memory\[342\]\[0\]
+ mod.u_cpu.rf_ram.memory\[343\]\[0\] _01826_ _01828_ _01840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_81_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_179_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_223_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_263_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07675__A1 _01934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07463_ _01569_ _01771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_223_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11471__A2 _05120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_222_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09202_ _03473_ _00029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__14780__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07394_ _01701_ _01702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07202__I _01509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_241_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07427__A1 _01493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09133_ _03363_ _03416_ _03426_ _03429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_176_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_191_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_191_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12971__A2 _06142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09064_ _03362_ _03363_ _03355_ _03364_ _03366_ _03367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_162_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_190_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15136__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08015_ _01665_ _02323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_135_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_200_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08927__A1 _02523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09129__I _03392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_190_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11782__I0 _05329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10585__I1 mod.u_cpu.rf_ram.memory\[428\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09966_ _04086_ _00183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__15286__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07872__I _01778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_265_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09727__I0 _03877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08917_ _02471_ _03216_ _03223_ _02491_ _03224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_103_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09897_ _04040_ _00160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11394__I _05031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08786__S0 _01673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08848_ mod.u_cpu.rf_ram.memory\[37\]\[1\] _03155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_57_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13287__I0 mod.u_arbiter.i_wb_cpu_rdt\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08779_ _01688_ _03078_ _03085_ _02291_ _03086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_27_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_232_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_245_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_150_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09799__I _03968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_168_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13987__A1 mod.u_arbiter.i_wb_cpu_rdt\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10810_ _03941_ _04668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_2847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_214_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11790_ _05338_ _00755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11837__I1 mod.u_cpu.rf_ram.memory\[228\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_198_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_214_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_214_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_198_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07666__A1 _01956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13039__I0 _06184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10741_ _04620_ _04621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_214_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_201_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_198_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13739__A1 _06713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_159_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13460_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[13\] _06531_ _06532_ _03569_ _06534_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_10672_ _04299_ _04575_ _04576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_179_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07418__A1 _01605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12411_ _02117_ _05758_ _05760_ _00954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_90_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_223_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_13391_ _06435_ _06486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_154_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13050__S _06201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07969__A2 _02268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15130_ _00983_ net3 mod.u_cpu.rf_ram.memory\[167\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10273__I0 _04298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_194_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08091__A1 _01823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12342_ _05494_ _05703_ _05714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_182_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10973__A1 _03663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08371__C _02677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14164__A1 _03298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_177_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15061_ _00915_ net3 mod.u_cpu.rf_ram.memory\[18\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_177_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12273_ _05666_ _05667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_49_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_218_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14503__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15629__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14012_ _03458_ _06964_ _06971_ mod.u_arbiter.i_wb_cpu_dbus_dat\[15\] _06972_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_11224_ _04795_ _04951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_153_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11773__I0 _05311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11155_ _04846_ _04905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_1_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07782__I _01661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10106_ _03835_ _04184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_49_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_255_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11086_ _04858_ _00531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_5451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_249_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11525__I0 _05147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14653__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14914_ _00768_ net3 mod.u_cpu.rf_ram.memory\[39\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10037_ _03992_ _04132_ _04134_ _04135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_114_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_209_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11150__A1 _04758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_237_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_224_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14845_ _00699_ net3 mod.u_cpu.rf_ram.memory\[265\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_4794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_208_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_184_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_251_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_217_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_205_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__15009__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__13978__A1 mod.u_arbiter.i_wb_cpu_dbus_dat\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14776_ _00630_ net3 mod.u_cpu.rf_ram.memory\[2\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_95_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11988_ _05448_ _05475_ _05476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_32_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08546__C _02852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_264_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_210_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07657__A1 _01963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13727_ _06417_ _06733_ _06321_ _06486_ _06734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_189_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12650__A1 _05293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10939_ _04719_ _04756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13024__I _06072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_204_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07752__S1 _01723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_176_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13658_ _06667_ _06669_ _06670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_158_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15159__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_220_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_12609_ _05887_ mod.u_cpu.rf_ram.memory\[153\]\[0\] _05897_ _05898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__11205__A2 _03986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12863__I _05786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12402__A1 _05300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13589_ _06615_ _01277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10264__I0 _04288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15328_ _01105_ net3 mod.u_cpu.rf_ram.memory\[409\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_185_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14155__A1 _06057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15259_ _00015_ net4 mod.u_arbiter.i_wb_cpu_rdt\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_160_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13902__A1 _03359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13902__B2 _06463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09582__A1 _03758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09820_ _03870_ _03966_ _03984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_154_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_247_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09751_ _03711_ _03779_ _03931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_67_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_228_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08702_ _02665_ _03000_ _03008_ _02852_ _03009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__08137__A2 _02425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09334__A1 _03554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09682_ _03876_ _00109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_41_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_251_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08633_ _02090_ _02939_ _02940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_230_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_215_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13643__B _06137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07440__S0 _01745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_214_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_227_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_208_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11819__I1 mod.u_cpu.rf_ram.memory\[230\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08564_ _01961_ _02867_ _02870_ _01972_ _02871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_74_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07515_ _01506_ _01823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08456__C _01698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08495_ _02041_ mod.u_cpu.rf_ram.memory\[332\]\[1\] _02801_ _02802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_211_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07446_ mod.u_cpu.rf_ram.memory\[421\]\[0\] _01754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_195_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_202_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_195_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12773__I _03734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07377_ _01680_ _01684_ _01685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_182_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14526__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_182_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09116_ _03414_ _03415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_182_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12944__A2 _06120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08073__A1 _02337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10955__A1 _04766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_237_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_164_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09047_ _03349_ _03296_ _03350_ _03250_ _03351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_159_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14676__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_237_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09949_ _04071_ mod.u_cpu.rf_ram.memory\[526\]\[1\] _04074_ _04076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_4002 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4013 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09325__A1 _03568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_219_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4024 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4035 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12960_ mod.u_arbiter.i_wb_cpu_ack _03399_ _06136_ _06137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_4046 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_161_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12180__I0 _05583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4057 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4068 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11911_ _05422_ _05423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_161_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4079 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07887__A1 _02188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_261_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_218_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12891_ _06083_ _01111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_166_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_233_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14630_ _00484_ net3 mod.u_cpu.rf_ram.memory\[372\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_45_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11842_ _05373_ _05374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1910 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1921 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1932 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_207_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07639__A1 _01934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1943 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14561_ _00415_ net3 mod.u_cpu.rf_ram.memory\[407\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_220_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11773_ _05311_ mod.u_cpu.rf_ram.memory\[236\]\[0\] _05326_ _05327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_1954 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15301__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_207_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1965 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1976 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08300__A2 _02598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13512_ _06567_ _01248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_10724_ _04184_ _04574_ _04610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1987 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14492_ _00346_ net3 mod.u_cpu.rf_ram.memory\[441\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1998 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_202_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13443_ _06523_ _01223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_10655_ _04560_ mod.u_cpu.rf_ram.memory\[417\]\[1\] _04562_ _04564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_155_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07777__I _02084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08064__A1 _02302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15451__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13374_ _06374_ _06470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_142_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_194_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10586_ _04517_ _00372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_182_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09800__A2 _03969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15113_ _00002_ net3 mod.u_cpu.cpu.alu.i_rs1 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_86_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12325_ _05692_ mod.u_cpu.rf_ram.memory\[179\]\[1\] _05700_ _05702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_154_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07811__A1 _02115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15044_ _00898_ net3 mod.u_cpu.rf_ram.memory\[109\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_114_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12256_ _05655_ _00904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_142_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_190_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11207_ _04940_ _00570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08367__A2 _02673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12187_ _05608_ _00882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_96_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_229_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11138_ _04749_ _04887_ _04894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_96_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09316__A1 _03563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_237_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11069_ _04846_ _04847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_5281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xtiny_user_project_140 la_data_out[58] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_76_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xtiny_user_project_151 wbs_dat_o[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_114_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xtiny_user_project_162 wbs_dat_o[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_225_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_237_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_149_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_173 wbs_dat_o[23] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__10579__S _04512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_209_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14828_ _00682_ net3 mod.u_cpu.rf_ram.memory\[273\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_91_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_52_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14759_ _00613_ net3 mod.u_cpu.rf_ram.memory\[308\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__13820__B1 _06466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_264_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_177_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_225_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07300_ _01510_ _01608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_60_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14549__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08280_ mod.u_cpu.rf_ram.memory\[461\]\[1\] _02587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_149_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07231_ _01538_ _01539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_20_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__12593__I _05694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_177_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_192_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07687__I _01762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07162_ _01470_ _01471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_121_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11985__I0 _05464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14699__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13351__A2 _06390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11362__A1 _05047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09803_ _03964_ mod.u_cpu.rf_ram.memory\[547\]\[1\] _03970_ _03972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_8_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_219_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07995_ _01862_ _02303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_228_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09734_ _03917_ _03918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_95_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07869__A1 _02157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09665_ _03863_ _00105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_67_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_243_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15324__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_215_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08616_ _02916_ _02918_ _02920_ _02922_ _01658_ _02923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_82_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09596_ _03809_ _03810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_199_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_231_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_243_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_202_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08547_ _02841_ _02843_ _01891_ _02853_ _02854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__12614__A1 _05283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_196_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08294__A1 _02585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15474__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13820__C _06776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08478_ _01875_ mod.u_cpu.rf_ram.memory\[366\]\[1\] _02784_ _02030_ _02785_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_196_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07429_ _01486_ _01736_ _01737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12217__I1 mod.u_cpu.rf_ram.memory\[198\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_183_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08046__A1 _02266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10440_ _04410_ mod.u_cpu.rf_ram.memory\[452\]\[1\] _04417_ _04419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_136_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08597__A2 mod.u_cpu.rf_ram.memory\[260\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10371_ _04363_ mod.u_cpu.rf_ram.memory\[463\]\[1\] _04370_ _04372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_87_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12110_ _05367_ _05543_ _05556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_124_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13090_ _06217_ mod.u_cpu.rf_ram.memory\[103\]\[1\] _06227_ _06229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_156_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13878__B1 _06866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12041_ _05510_ _00834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13342__A2 _06390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_215_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_215_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_213_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13992_ _06955_ _06956_ _01339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_77_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09849__A2 _03996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_248_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_12943_ _05784_ _03458_ _06119_ _06120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_3120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_234_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10399__S _04390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_234_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08521__A2 mod.u_cpu.rf_ram.memory\[340\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_206_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12874_ _03923_ _06072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_234_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11825_ _05361_ _00767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_14613_ _00467_ net3 mod.u_cpu.rf_ram.memory\[381\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_15593_ _01364_ net3 mod.u_cpu.rf_ram.memory\[299\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_92_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_221_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_199_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14544_ _00398_ net3 mod.u_cpu.rf_ram.memory\[415\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11756_ _05304_ mod.u_cpu.rf_ram.memory\[238\]\[1\] _05313_ _05315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_1784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_222_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__13730__C _06640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_201_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10092__A1 _04172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_187_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10707_ _04574_ _04599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_105_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14841__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_187_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14475_ _00329_ net3 mod.u_cpu.rf_ram.memory\[450\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11687_ _05267_ _00723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_197_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_146_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08037__A1 _01493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13426_ _06512_ _06513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_10638_ _04537_ mod.u_cpu.rf_ram.memory\[420\]\[1\] _04551_ _04553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__13030__A1 _03904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07300__I _01510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13357_ _06449_ _06451_ _06452_ _06453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_154_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10569_ _04505_ _00367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_182_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10395__A2 _03807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__14991__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_182_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12308_ _04873_ _05686_ _05690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_115_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13288_ _06377_ mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat\[2\] _06386_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_114_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15027_ _00881_ net3 mod.u_cpu.rf_ram.memory\[204\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12239_ mod.u_cpu.rf_ram.memory\[109\]\[1\] _05617_ _05641_ _05644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_142_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_256_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15347__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08760__A2 _03059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14133__I1 mod.u_cpu.rf_ram.memory\[115\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07780_ _02083_ _02087_ _02088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_111_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12144__I0 _05566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput4 io_in[8] net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_12
Xtiny_user_project_90 la_data_out[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_225_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12695__I1 _05950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12844__A1 _05788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_266_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_266_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_252_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09450_ mod.u_arbiter.i_wb_cpu_ibus_adr\[0\] mod.u_cpu.cpu.ctrl.pc_plus_offset_cy_r
+ _03265_ _03678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_188_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14371__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__15497__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_266_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08401_ _02692_ mod.u_cpu.rf_ram.memory\[438\]\[1\] _02707_ _01981_ _02708_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_91_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_197_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09381_ _03618_ _03619_ _03620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_80_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_221_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08332_ mod.u_cpu.rf_ram.memory\[503\]\[1\] _02639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__10458__I0 _04430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_178_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08276__A1 _01464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_162_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_177_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08263_ _02523_ _02562_ _02570_ _02469_ _02571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__13212__I _06318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07214_ _01520_ _01521_ _01522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08194_ _02500_ _02501_ _02502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07210__I _01515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07145_ mod.u_cpu.cpu.decode.op26 _01453_ _01454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_238_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_134_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07251__A2 mod.u_cpu.rf_ram.memory\[476\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_161_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11335__A1 _04196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_259_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_248_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10933__I1 mod.u_cpu.rf_ram.memory\[372\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08751__A2 _03057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13088__A1 _06032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07978_ _02129_ mod.u_cpu.rf_ram.memory\[100\]\[0\] _02285_ _02286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_59_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12135__I0 _05559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14714__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07880__I _01582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09717_ _03904_ _03905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07813__C _02120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_228_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_83_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09648_ _03849_ _03850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_216_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_216_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_231_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09801__S _03970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14864__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09579_ _03745_ _03786_ _03795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12438__I1 mod.u_cpu.rf_ram.memory\[172\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10947__S _04760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_203_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_167_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11610_ _05119_ _05214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10449__I0 _04423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08267__A1 _02546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_230_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_212_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12063__A2 _03771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_12590_ _05884_ _01009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_168_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_212_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08644__C _01771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11541_ _05159_ mod.u_cpu.rf_ram.memory\[276\]\[0\] _05168_ _05169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_196_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_212_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07865__I1 mod.u_cpu.rf_ram.memory\[201\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11810__A2 _03866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_211_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14260_ _00114_ net3 mod.u_cpu.rf_ram.memory\[557\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08019__A1 _02298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11472_ _05022_ _05121_ _05122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__13012__A1 _03837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_221_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07490__A2 mod.u_cpu.rf_ram.memory\[438\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_183_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_13211_ _06317_ _06318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_10423_ _04308_ _04407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08114__S1 _02350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14191_ _07091_ _01403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12961__I _06137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13142_ _06261_ _01184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_139_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10354_ _03865_ _04360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__14244__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13073_ _06217_ mod.u_cpu.rf_ram.memory\[81\]\[1\] _06215_ _06218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_151_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10285_ _04313_ mod.u_cpu.rf_ram.memory\[477\]\[1\] _04310_ _04314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_3_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12024_ _05498_ mod.u_cpu.rf_ram.memory\[58\]\[0\] _05499_ _05500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__13866__A3 _06858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07625__S0 _01802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11877__A2 _05398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_238_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14394__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_266_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_265_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__12126__I0 _05566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13725__C _06713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07790__I _01637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_254_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_266_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_219_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_207_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11629__A2 _05210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12826__A1 _06032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07723__C _02030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13975_ mod.u_arbiter.i_wb_cpu_dbus_dat\[7\] _06943_ _06944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_81_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_207_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11018__S _04809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_234_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09542__I1 mod.u_cpu.rf_ram.memory\[574\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10688__I0 _04579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_234_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12926_ _06106_ _01123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_18_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_261_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15645_ _01416_ net3 mod.u_cpu.rf_ram.memory\[249\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_222_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12857_ _01464_ mod.u_cpu.rf_ram.regzero _06059_ _01101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XTAP_2271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_226_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11808_ _05350_ mod.u_cpu.rf_ram.memory\[231\]\[1\] _05347_ _05351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_61_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15576_ _01347_ net3 mod.u_arbiter.i_wb_cpu_dbus_dat\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12788_ _03974_ _06011_ _06015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_187_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09510__I _03734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10065__A1 _03791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08554__C _01952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11739_ _05289_ mod.u_cpu.rf_ram.memory\[240\]\[0\] _05302_ _05303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_175_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14527_ _00381_ net3 mod.u_cpu.rf_ram.memory\[424\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_230_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_14458_ _00312_ net3 mod.u_cpu.rf_ram.memory\[458\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07481__A2 _01772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_179_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12871__I _06018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13409_ _06501_ _01211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_122_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_14389_ _00243_ net3 mod.u_cpu.rf_ram.memory\[493\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_143_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10368__A2 _04335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10612__I0 _04523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11487__I _05132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08950_ _03254_ _03255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_143_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08997__S mod.u_cpu.rf_ram_if.rtrig1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14737__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12365__I0 _05729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07901_ _02091_ _02209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_142_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08881_ mod.u_cpu.rf_ram.memory\[573\]\[1\] _03188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_155_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11868__A2 _05388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_257_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07832_ _02135_ mod.u_cpu.rf_ram.memory\[166\]\[0\] _02138_ _02139_ _02140_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_57_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12312__S _05690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12117__I0 _05559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08729__C _01702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07763_ _01746_ _02071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__14887__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07633__C _01783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_186_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09502_ _03723_ _03727_ _03728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_253_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_225_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08497__A1 _02672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07694_ mod.u_cpu.rf_ram.memory\[287\]\[0\] _02002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__14019__B1 _06971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13490__A1 _03616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11340__I1 mod.u_cpu.rf_ram.memory\[30\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09433_ mod.u_cpu.cpu.immdec.imm11_7\[2\] _03664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08592__S1 _01932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_266_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__10767__S _04638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_213_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_240_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_212_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08249__A1 _02542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09364_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[22\] _03605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12045__A2 _05512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_244_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08315_ _02225_ _02621_ _02622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_177_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09295_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[11\] _03547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_166_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08246_ _02550_ mod.u_cpu.rf_ram.memory\[526\]\[0\] _02553_ _02515_ _02554_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_36_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14267__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15512__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_180_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08177_ mod.u_cpu.rf_ram.memory\[559\]\[0\] _02485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_153_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_192_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07128_ _01433_ _01434_ _01436_ _01437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__08421__A1 _02244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11397__I _05045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08811__I3 mod.u_cpu.rf_ram.memory\[3\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08972__A2 _03270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10070_ _04158_ _00215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13826__B _06490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_247_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_236_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__12108__I0 _05550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_229_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_210_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12808__A1 _02234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_216_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13760_ mod.u_cpu.cpu.immdec.imm31 _03274_ _06764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_28_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08488__A1 _02668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10972_ _04778_ _00497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08032__S0 _01857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_210_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_243_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_216_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12711_ _05965_ _01049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_253_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_13691_ mod.u_cpu.cpu.immdec.imm19_12_20\[3\] _06678_ _06701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_245_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_188_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15042__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12642_ _05372_ _05919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_15430_ _01205_ net3 mod.u_cpu.rf_ram.memory\[95\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_169_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_231_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13233__B2 _06339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_197_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15361_ _01136_ net3 mod.u_cpu.rf_ram.memory\[86\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__13784__A2 _06783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12573_ _05709_ _05873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_157_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_196_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_200_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11524_ _05157_ _00670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_141_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14312_ _00166_ net3 mod.u_cpu.rf_ram.memory\[531\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_15292_ _00051_ net4 mod.u_scanchain_local.module_data_in\[49\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_183_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08660__A1 _02656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_183_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15192__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14243_ _00097_ net3 mod.u_cpu.rf_ram.memory\[566\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_144_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11455_ _05109_ _00649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_172_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10406_ _03924_ _04396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_125_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14174_ _03928_ _07081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08412__A1 _02654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11386_ _04817_ _05063_ _05064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_178_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13125_ _06251_ _01177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_10337_ _04189_ _04327_ _04349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_113_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11100__I _03795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13056_ _06207_ _01152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_10268_ _03721_ _04133_ _04300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_65_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12007_ _05488_ _05486_ _05489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_117_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10199_ _04249_ mod.u_cpu.rf_ram.memory\[48\]\[0\] _04252_ _04253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07923__B1 _02229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_235_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08479__A1 _01997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13958_ _03441_ _05793_ _06930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_47_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12275__A2 _05668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_222_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12909_ _06095_ _01117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_228_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_222_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13889_ _06868_ _06836_ _06872_ _06880_ _01312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_50_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_222_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15628_ _01399_ net3 mod.u_cpu.rf_ram.memory\[8\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_146_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2090 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_222_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09240__I _03500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_203_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__15535__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10386__I _03928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_187_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15559_ _01330_ net3 mod.u_arbiter.i_wb_cpu_dbus_dat\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_188_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_187_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11786__A1 _05334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08100_ _02406_ _02407_ _02408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_175_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10589__A2 _04507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09080_ _03378_ _03381_ _03382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_238_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_135_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08031_ _02090_ _02338_ _02339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09396__B _03493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_200_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_174_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11389__I1 _05065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07206__A2 mod.u_cpu.rf_ram.memory\[452\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10061__I1 mod.u_cpu.rf_ram.memory\[508\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09982_ _04096_ mod.u_cpu.rf_ram.memory\[520\]\[0\] _04097_ _04098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_116_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08933_ _02551_ _03239_ _03240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_83_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_233_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11010__I0 _04803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09903__A1 _04044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12042__S _05509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08864_ _02456_ mod.u_cpu.rf_ram.memory\[548\]\[1\] _03170_ _03171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_97_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_229_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_170_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_218_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07815_ _01670_ _02108_ _02121_ _02122_ _02123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_96_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08795_ _02465_ _03098_ _03101_ _02660_ _03102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_211_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07746_ _01569_ _02054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__15065__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_225_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_203_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12510__I0 _05827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09131__A2 _03387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07677_ mod.u_cpu.rf_ram.memory\[279\]\[0\] _01985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__11680__I _05253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_164_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_241_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_198_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09416_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[29\] mod.u_cpu.cpu.ctrl.o_ibus_adr\[28\] _03635_
+ _03632_ _03650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_53_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07693__A2 mod.u_cpu.rf_ram.memory\[284\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10029__A1 _03986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09150__I _03417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_209_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_201_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09347_ _03436_ mod.u_scanchain_local.module_data_in\[55\] _03402_ mod.u_arbiter.i_wb_cpu_dbus_adr\[18\]
+ _03592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_205_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_197_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13766__A2 _06753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_240_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13601__S _06621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14902__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09278_ _03525_ _03532_ _03533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_201_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_194_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08229_ _01747_ _02537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13400__I _06434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_193_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11240_ _04963_ _00580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_165_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11171_ _04879_ _04916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12016__I _03827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12329__I0 _05696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10122_ _04195_ _04196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_122_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_5600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_251_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14930_ _00784_ net3 mod.u_cpu.rf_ram.memory\[227\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09745__I1 _03925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10053_ _03738_ _04147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_5644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_209_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4910 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15408__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4921 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_209_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_76_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4932 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08369__C _01687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_180_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4943 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14861_ _00715_ net3 mod.u_cpu.rf_ram.memory\[258\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_169_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4954 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_180_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13829__I0 mod.u_arbiter.i_wb_cpu_rdt\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_264_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4965 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4976 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_180_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4987 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13812_ _06482_ _06772_ _06812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_29_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_217_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4998 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14792_ _00646_ net3 mod.u_cpu.rf_ram.memory\[291\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_113_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_249_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_217_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10268__A1 _03721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_232_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_204_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13743_ _06678_ _06456_ _06742_ _06748_ _06749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
X_10955_ _04766_ _04759_ _04767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__15558__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14432__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_204_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13674_ _06304_ _06370_ _06682_ _06661_ _06684_ _06306_ _06685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_143_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10886_ _04720_ mod.u_cpu.rf_ram.memory\[380\]\[1\] _04717_ _04721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_71_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15413_ _01188_ net3 mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_12625_ _05908_ _01020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_197_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_185_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__14582__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10815__I0 _04666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15344_ _01119_ net3 mod.u_cpu.rf_ram.memory\[399\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08633__A1 _02090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12556_ _05858_ mod.u_cpu.rf_ram.memory\[162\]\[1\] _05860_ _05862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_223_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_200_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_184_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11507_ _05146_ _00664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_185_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08832__C _02363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13509__A2 _03302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_200_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10291__I1 mod.u_cpu.rf_ram.memory\[476\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15275_ _00033_ net4 mod.u_arbiter.i_wb_cpu_rdt\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_8_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__12980__A3 _06151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12487_ _05813_ mod.u_cpu.rf_ram.memory\[171\]\[0\] _05817_ _05818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_176_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14226_ _00080_ net3 mod.u_cpu.rf_ram.memory\[574\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__14182__A2 _05124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11438_ _05096_ mod.u_cpu.rf_ram.memory\[292\]\[0\] _05097_ _05098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_208_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_171_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_256_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_153_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11966__S _05459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08936__A2 _03235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14157_ _06056_ mod.u_cpu.cpu.state.o_cnt_r\[2\] _07069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_11369_ _05046_ mod.u_cpu.rf_ram.memory\[304\]\[0\] _05052_ _05053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_28_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_193_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08492__S0 _01920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_217_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11940__A1 _05443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13108_ mod.u_cpu.rf_ram.memory\[101\]\[1\] _06221_ _06239_ _06241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_14088_ _03836_ _05279_ _07025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_98_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13039_ _06184_ mod.u_cpu.rf_ram.memory\[83\]\[1\] _06194_ _06196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__15088__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_230_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09235__I _03495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11543__I1 mod.u_cpu.rf_ram.memory\[276\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_67_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_227_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_227_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07600_ _01745_ mod.u_cpu.rf_ram.memory\[358\]\[0\] _01907_ _01882_ _01908_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_93_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_254_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_208_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08580_ _01998_ mod.u_cpu.rf_ram.memory\[284\]\[1\] _02886_ _02887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_82_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_207_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07531_ mod.u_cpu.rf_ram.memory\[324\]\[0\] mod.u_cpu.rf_ram.memory\[325\]\[0\] mod.u_cpu.rf_ram.memory\[326\]\[0\]
+ mod.u_cpu.rf_ram.memory\[327\]\[0\] _01837_ _01838_ _01839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__07911__C _02218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_223_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11206__S _04939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_223_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_228_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_223_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_179_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07514__I3 mod.u_cpu.rf_ram.memory\[335\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07462_ _01741_ _01770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__14925__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07675__A2 _01982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08872__A1 _02479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_250_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09201_ mod.u_arbiter.i_wb_cpu_rdt\[26\] mod.u_arbiter.i_wb_cpu_dbus_dat\[23\] _03469_
+ _03473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_179_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07393_ _01700_ _01701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_72_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_210_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_241_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_188_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09416__A3 _03635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09132_ mod.u_arbiter.i_wb_cpu_rdt\[2\] _03428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_249_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07427__A2 _01724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08624__A1 _02074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_176_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10431__A1 _04412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09063_ _03354_ _03365_ _03366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__12037__S _05506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12559__I0 _05855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_194_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08014_ _02293_ _02312_ _02320_ _02321_ _02322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_191_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_239_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08927__A2 _03226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14305__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09965_ _04071_ mod.u_cpu.rf_ram.memory\[523\]\[1\] _04084_ _04086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_258_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09727__I1 mod.u_cpu.rf_ram.memory\[555\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08916_ _02545_ _03219_ _03222_ _02489_ _03223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__14051__I _06914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09896_ _04023_ mod.u_cpu.rf_ram.memory\[534\]\[0\] _04039_ _04040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_134_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_170_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_170_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08847_ mod.u_cpu.rf_ram.memory\[32\]\[1\] mod.u_cpu.rf_ram.memory\[33\]\[1\] mod.u_cpu.rf_ram.memory\[34\]\[1\]
+ mod.u_cpu.rf_ram.memory\[35\]\[1\] _01647_ _01732_ _03154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_3505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14455__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08786__S1 _01855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_257_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13890__I _06704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08778_ _02325_ _03081_ _03084_ _01717_ _03085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_72_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_233_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13287__I1 mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_226_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07729_ _01471_ _01913_ _02036_ _02037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__08917__C _02491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_198_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13987__A2 _06952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_226_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_214_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_198_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_207_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11998__A1 _05448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10740_ _03737_ _04620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_214_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07666__A2 _01959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08863__A1 _02472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_240_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13739__A2 _06744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10671_ _04574_ _04575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_198_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_201_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_12410_ _05759_ _05758_ _05760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_90_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13390_ _05784_ mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat\[10\] _06484_ _06485_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__08615__A1 _02057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12411__A2 _05758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12341_ _05695_ _05713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_182_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10273__I1 mod.u_cpu.rf_ram.memory\[478\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_216_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_194_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10973__A2 _04223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15060_ _00914_ net3 mod.u_cpu.rf_ram.memory\[18\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_138_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12272_ _03755_ _05371_ _05666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_181_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_257_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14011_ _06970_ _06971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11222__I0 _04938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11223_ _04950_ _00576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_175_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10025__I1 _03925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13911__A2 _06890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09040__A1 mod.u_cpu.cpu.state.o_cnt_r\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15230__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11773__I1 mod.u_cpu.rf_ram.memory\[236\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11154_ _04904_ _00553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_122_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10105_ _04183_ _00225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_95_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11085_ _04841_ mod.u_cpu.rf_ram.memory\[34\]\[1\] _04856_ _04858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_27_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13675__A1 _06431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_248_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_209_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11525__I1 mod.u_cpu.rf_ram.memory\[27\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_209_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14913_ _00767_ net3 mod.u_cpu.rf_ram.memory\[22\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10036_ _04133_ _04134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_5474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15380__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_236_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14844_ _00698_ net3 mod.u_cpu.rf_ram.memory\[265\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_4773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14948__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_263_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10929__I _03841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_205_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14775_ _00629_ net3 mod.u_cpu.rf_ram.memory\[300\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11987_ _03834_ _04068_ _05475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_147_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_205_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13305__I _06402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_95_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_260_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_13726_ _06438_ _06711_ _06733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_44_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_220_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07657__A2 _01964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08854__A1 _02063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10938_ _04755_ _00486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_232_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13657_ _06361_ _06668_ _06669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_10869_ _04708_ _04709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_34_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12789__I0 _06010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_176_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08606__A1 _01470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_12608_ _05896_ _05882_ _05897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__12402__A2 _05726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13588_ mod.u_arbiter.i_wb_cpu_dbus_adr\[26\] mod.u_arbiter.i_wb_cpu_dbus_adr\[27\]
+ _06614_ _06615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_200_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_191_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10413__A1 _04255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_185_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15327_ _01104_ net3 mod.u_cpu.rf_ram.memory\[409\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_117_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12539_ mod.u_cpu.rf_ram.memory\[165\]\[1\] _05765_ _05849_ _05851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_121_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__14328__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15258_ _00014_ net4 mod.u_arbiter.i_wb_cpu_rdt\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12166__A1 _04379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11213__I0 _04936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14209_ _02023_ _07100_ _07101_ _01412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_144_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15189_ _01042_ net3 mod.u_cpu.rf_ram.memory\[77\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_99_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_99_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09582__A2 _03797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14478__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07593__A1 _01852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09750_ _03930_ _00123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_234_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__12713__I0 _05966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08701_ _02063_ _03004_ _03007_ _01669_ _03008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_95_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09681_ _03862_ mod.u_cpu.rf_ram.memory\[560\]\[1\] _03874_ _03876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_239_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07345__A1 _01632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08632_ mod.u_cpu.rf_ram.memory\[184\]\[1\] mod.u_cpu.rf_ram.memory\[185\]\[1\] mod.u_cpu.rf_ram.memory\[186\]\[1\]
+ mod.u_cpu.rf_ram.memory\[187\]\[1\] _02092_ _02098_ _02939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_54_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12320__S _05697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_255_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07440__S1 _01747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_215_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08563_ _01697_ mod.u_cpu.rf_ram.memory\[310\]\[1\] _02869_ _01970_ _02870_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_70_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09098__A1 _03398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07514_ mod.u_cpu.rf_ram.memory\[332\]\[0\] mod.u_cpu.rf_ram.memory\[333\]\[0\] mod.u_cpu.rf_ram.memory\[334\]\[0\]
+ mod.u_cpu.rf_ram.memory\[335\]\[0\] _01819_ _01821_ _01822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_23_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_223_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14218__I0 _03699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08494_ _01729_ _02800_ _02801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_35_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_251_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_222_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07445_ _01752_ _01753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_167_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10652__A1 _04285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15103__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_211_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_183_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07376_ mod.u_cpu.rf_ram.memory\[392\]\[0\] mod.u_cpu.rf_ram.memory\[393\]\[0\] mod.u_cpu.rf_ram.memory\[394\]\[0\]
+ mod.u_cpu.rf_ram.memory\[395\]\[0\] _01682_ _01683_ _01684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_176_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_210_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09115_ _03413_ _03414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_148_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_198_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08073__A2 _02346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15253__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10955__A2 _04759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_191_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_136_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09046_ _03349_ _03316_ _03350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_198_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08044__I _01882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_191_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_150_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08979__I mod.u_cpu.cpu.state.init_done vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11904__A1 _05417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07883__I _02190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_35 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09948_ _04075_ _00176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_4003 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4014 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4025 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4036 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_161_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09879_ _04028_ _00154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_57_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4047 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12180__I1 mod.u_cpu.rf_ram.memory\[204\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4058 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_218_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4069 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11910_ _05421_ _05422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07887__A2 _02189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10191__I0 _04245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12890_ _06070_ mod.u_cpu.rf_ram.memory\[89\]\[1\] _06081_ _06083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_72_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11841_ _05372_ _05373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09089__A1 mod.u_cpu.cpu.state.o_cnt_r\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1900 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1911 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1922 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_242_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1933 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11772_ _05325_ _05301_ _05326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_202_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14560_ _00414_ net3 mod.u_cpu.rf_ram.memory\[407\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08219__I _02526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1944 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_214_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1955 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1966 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_186_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10723_ _04609_ _00417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1977 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13511_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[31\] _06557_ _06558_ _06566_ _06567_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_158_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_241_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_198_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14491_ _00345_ net3 mod.u_cpu.rf_ram.memory\[442\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1988 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1999 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__13188__A3 _06281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10654_ _04563_ _00394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_16_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_13442_ _03524_ _06519_ _06520_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[7\] _06523_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__12396__A1 _04700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11443__I0 _05096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13373_ _06468_ _06403_ _06469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08064__A2 mod.u_cpu.rf_ram.memory\[76\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10585_ _04506_ mod.u_cpu.rf_ram.memory\[428\]\[0\] _04516_ _04517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09261__A1 _03506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15112_ _00966_ net3 mod.u_cpu.raddr\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12324_ _05701_ _00926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_177_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12148__A1 _05581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14620__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12255_ _05645_ mod.u_cpu.rf_ram.memory\[194\]\[0\] _05654_ _05655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_15043_ _00897_ net3 mod.u_cpu.rf_ram.memory\[197\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_126_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09013__A1 _01431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11206_ _04938_ mod.u_cpu.rf_ram.memory\[32\]\[0\] _04939_ _04940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_79_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12186_ _05605_ mod.u_cpu.rf_ram.memory\[203\]\[0\] _05607_ _05608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07575__A1 _01879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_253_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_150_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11137_ _04893_ _00547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_150_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13648__A1 _06289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14770__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_249_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11068_ _04300_ _04701_ _04846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_231_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_95_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xtiny_user_project_130 la_data_out[48] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_5282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xtiny_user_project_141 la_data_out[59] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__13236__S _06341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_49_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10019_ _04117_ mod.u_cpu.rf_ram.memory\[514\]\[0\] _04122_ _04123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xtiny_user_project_152 wbs_dat_o[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_110_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_163 wbs_dat_o[13] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_36_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_225_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07878__A2 _02173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtiny_user_project_174 wbs_dat_o[24] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__10182__I0 _04217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09513__I _03695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_251_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14827_ _00681_ net3 mod.u_cpu.rf_ram.memory\[274\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__15126__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07461__C _01768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13035__I _05396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14758_ _00612_ net3 mod.u_cpu.rf_ram.memory\[308\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08827__A1 _02316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13820__A1 _06311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_233_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13820__B2 _06372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_204_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13709_ _06380_ _06448_ _06717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_149_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_220_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14689_ _00543_ net3 mod.u_cpu.rf_ram.memory\[343\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_220_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15276__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07230_ _01537_ _01538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_81_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_220_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07161_ _01463_ mod.u_cpu.cpu.immdec.imm19_12_20\[7\] _01467_ mod.u_cpu.cpu.immdec.imm24_20\[3\]
+ _01470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_173_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_146_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11985__I1 mod.u_cpu.rf_ram.memory\[216\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_246_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_145_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08438__S0 _02020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13887__A1 _06823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13887__B2 _06423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09802_ _03971_ _00134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_119_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07994_ _02134_ _02302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_140_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_228_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07208__I _01515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09733_ _03711_ _03745_ _03917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_228_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07318__A1 _01578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_228_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09664_ _03862_ mod.u_cpu.rf_ram.memory\[562\]\[1\] _03860_ _03863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08610__S0 _02085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_228_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08467__C _01867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_227_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08615_ _02057_ _02921_ _01632_ _02922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09595_ _03808_ _03809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_167_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_167_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13111__I0 _06230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_224_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_208_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08818__A1 _02302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08546_ _02196_ _02844_ _02851_ _02852_ _02853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__15619__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09866__I0 _04018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_211_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_196_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10625__A1 _04262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_223_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11673__I0 _05250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08477_ _02027_ _02783_ _02784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_126_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08294__A2 mod.u_cpu.rf_ram.memory\[452\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07428_ _01446_ _01721_ _01735_ _01736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_211_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_17_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_196_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_149_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_206_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__14643__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07359_ mod.u_cpu.rf_ram.memory\[384\]\[0\] mod.u_cpu.rf_ram.memory\[385\]\[0\] mod.u_cpu.rf_ram.memory\[386\]\[0\]
+ mod.u_cpu.rf_ram.memory\[387\]\[0\] _01664_ _01666_ _01667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__08046__A2 _02353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10370_ _01546_ _04370_ _04371_ _00302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_191_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09029_ _03302_ _03333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_3_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14793__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12040_ _05498_ mod.u_cpu.rf_ram.memory\[60\]\[0\] _05509_ _05510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12925__I0 _06105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_176_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_254_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15149__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13991_ _03449_ _06952_ _06947_ mod.u_arbiter.i_wb_cpu_dbus_dat\[10\] _06956_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_120_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_213_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08658__B _01738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_219_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12942_ _03500_ mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat\[15\] _06119_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_3121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_233_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10864__A1 _04611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12873_ _06071_ _01105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_215_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15299__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14612_ _00466_ net3 mod.u_cpu.rf_ram.memory\[381\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11824_ _05350_ mod.u_cpu.rf_ram.memory\[22\]\[1\] _05359_ _05361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08809__A1 _01483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15592_ _01363_ net3 mod.u_cpu.rf_ram.memory\[299\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__13802__A1 _06418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09857__I0 _03999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_202_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13802__B2 _06443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11664__I0 _05250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_187_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14543_ _00397_ net3 mod.u_cpu.rf_ram.memory\[416\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11755_ _05314_ _00744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_199_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_187_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07788__I _01686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_202_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_202_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10706_ _04522_ _04598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_14474_ _00328_ net3 mod.u_cpu.rf_ram.memory\[450\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_105_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11686_ _05250_ mod.u_cpu.rf_ram.memory\[255\]\[1\] _05264_ _05267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_202_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12369__A1 _05732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_174_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13425_ net5 _03677_ _06512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_155_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10637_ _04552_ _00388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_167_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13030__A2 _06092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13356_ _06426_ _06452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_10568_ _04498_ mod.u_cpu.rf_ram.memory\[431\]\[1\] _04503_ _04505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_182_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_220_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10942__I _03857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12307_ _05689_ _00921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_114_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13869__A1 _06694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13287_ mod.u_arbiter.i_wb_cpu_rdt\[3\] mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat\[3\]
+ _06377_ _06385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_10499_ _04450_ mod.u_cpu.rf_ram.memory\[443\]\[1\] _04458_ _04460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_170_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09508__I _03732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15026_ _00880_ net3 mod.u_cpu.rf_ram.memory\[204\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_216_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_12238_ _02299_ _05641_ _05643_ _00898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07456__C _01763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_190_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12541__A1 _05367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12169_ _02176_ _05595_ _05596_ _00876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_29_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_190_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_80 io_out[36] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xinput5 io_in[9] net5 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xtiny_user_project_91 la_data_out[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_5090 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14516__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12844__A2 _05803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_237_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_209_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_264_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_225_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_227_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_225_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08400_ _01709_ _02706_ _02707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_206_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09380_ _03616_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[23\] mod.u_cpu.cpu.ctrl.o_ibus_adr\[22\]
+ _03619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_52_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13921__C _06481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_252_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_196_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08331_ _01537_ _02638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__11655__I0 _05243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14666__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10458__I1 mod.u_cpu.rf_ram.memory\[44\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_178_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08276__A2 _01465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08262_ _02525_ _02565_ _02569_ _02539_ _02570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_60_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_221_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_178_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07213_ mod.u_cpu.rf_ram.memory\[455\]\[0\] _01521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_220_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_192_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08193_ mod.u_cpu.rf_ram.memory\[575\]\[0\] _02501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__08028__A2 _02311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_257_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07144_ mod.u_cpu.cpu.decode.co_ebreak _01453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_119_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09776__A2 _03951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07787__A1 _02090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07331__S0 _01636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07539__A1 _01836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11335__A2 _03752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12532__A1 _05642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_236_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13088__A2 _06227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07977_ _02130_ _02284_ _02285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_102_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11683__I _05132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09716_ _03903_ _03904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_132_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_262_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_256_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_216_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15441__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_216_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_215_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11894__I0 _05406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09647_ _03788_ _03848_ _03849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_16_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07711__A1 _01956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_204_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08992__I _03251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09578_ _03794_ _00087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09839__I0 _03999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_212_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_212_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08529_ _02148_ _02798_ _02835_ _02836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__10449__I1 mod.u_cpu.rf_ram.memory\[450\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_23_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15591__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_212_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11540_ _04749_ _05149_ _05168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11271__A1 _04983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_204_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_204_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11471_ _04700_ _05120_ _05121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_168_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13012__A2 _06080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13210_ _06309_ _06316_ _06317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10422_ _04406_ _00319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12071__I0 _05518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14190_ _07081_ mod.u_cpu.rf_ram.memory\[244\]\[1\] _07089_ _07091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_104_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08814__I1 _03118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_167_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_192_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13141_ mod.u_arbiter.i_wb_cpu_rdt\[22\] mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat\[6\]
+ _06258_ _06261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_137_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10353_ _04359_ _00297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_124_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13072_ _06104_ _06217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_10284_ _04266_ _04313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_2_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11326__A2 _05021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11794__S _05339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_183_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12023_ _05452_ _03810_ _05499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_105_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_254_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__13720__B1 _06725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_215_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07625__S1 _01932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14539__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08742__A3 _03048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12126__I1 mod.u_cpu.rf_ram.memory\[20\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_207_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_13974_ _06942_ _06943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10137__I0 _04193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12826__A2 _06040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_219_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_207_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14689__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12925_ _06105_ mod.u_cpu.rf_ram.memory\[379\]\[1\] _06102_ _06106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_246_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09998__I _04107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_207_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10002__I _03928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15644_ _01415_ net3 mod.u_cpu.rf_ram.memory\[259\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_73_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12856_ mod.u_cpu.rf_ram.rdata\[1\] _06059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_62_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_221_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_178_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_265_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11637__I0 _05222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11807_ _05328_ _05350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_2294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15575_ _01346_ net3 mod.u_arbiter.i_wb_cpu_dbus_dat\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09455__A1 _03349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08889__S0 _02457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12787_ _06014_ _01076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_30_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10065__A2 _04143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14526_ _00380_ net3 mod.u_cpu.rf_ram.memory\[424\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11738_ _05300_ _05301_ _05302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_203_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_202_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_174_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14457_ _00311_ net3 mod.u_cpu.rf_ram.memory\[45\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11669_ _05254_ _05255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__14200__A1 _06046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_13408_ _06351_ mod.u_cpu.rf_ram.memory\[91\]\[0\] _06500_ _06501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_190_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14388_ _00242_ net3 mod.u_cpu.rf_ram.memory\[493\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07313__S0 _01605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15314__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_196_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13339_ _06434_ _06435_ _06436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_115_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09238__I _03498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08142__I _02209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_233_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12514__A1 _05395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15009_ _00863_ net3 mod.u_cpu.rf_ram.memory\[20\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_07900_ _02196_ _02201_ _02206_ _02207_ _02208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_102_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08880_ mod.u_cpu.rf_ram.memory\[568\]\[1\] mod.u_cpu.rf_ram.memory\[569\]\[1\] mod.u_cpu.rf_ram.memory\[570\]\[1\]
+ mod.u_cpu.rf_ram.memory\[571\]\[1\] _02494_ _02451_ _03187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_116_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08813__S0 _02171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_256_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08194__A1 _02500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15464__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07831_ _01746_ _02139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_69_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_97_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__12599__I _05873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12117__I1 mod.u_cpu.rf_ram.memory\[210\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_244_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07762_ _01806_ _02070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_238_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_266_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09501_ _03726_ _03727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__10828__A1 _04272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07693_ _01998_ mod.u_cpu.rf_ram.memory\[284\]\[0\] _02000_ _02001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__14019__A1 mod.u_arbiter.i_wb_cpu_rdt\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13932__B _03279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08497__A2 _02803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11008__I _03931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09432_ _03662_ _03663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_92_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_198_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_266_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_80_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_197_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13778__B1 _06779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09363_ _03489_ _03603_ _03604_ _00062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__08249__A2 _02544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09446__A1 _03371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13223__I _06329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08314_ mod.u_cpu.rf_ram.memory\[469\]\[1\] _02621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_162_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09294_ _03488_ _03546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_205_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10300__I0 _04298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07221__I _01528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_205_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_193_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11879__S _05398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08245_ _02551_ _02552_ _02553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_165_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_203_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_197_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08761__B _02149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_197_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08176_ _01745_ _02484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_14_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_238_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08480__C _02007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07127_ _01435_ _01420_ _01423_ _01436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_133_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_248_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_212_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14831__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07932__A1 _02155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12302__I _05667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12808__A2 _06027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_263_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_228_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08327__I3 mod.u_cpu.rf_ram.memory\[499\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10971_ _04772_ mod.u_cpu.rf_ram.memory\[366\]\[1\] _04776_ _04778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10958__S _04767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08032__S1 _02054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08732__I0 mod.u_cpu.rf_ram.memory\[248\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_210_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12710_ _05963_ mod.u_cpu.rf_ram.memory\[7\]\[0\] _05964_ _05965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_71_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11492__A1 _04859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_216_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13690_ _06693_ _06463_ _06699_ _06409_ _06700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_216_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_203_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__14981__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11619__I0 _05208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08655__C _02143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07791__S0 _02092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12641_ _05886_ _05918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_31_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09437__A1 _03289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_246_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_71_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11244__A1 _04965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15360_ _01135_ net3 mod.u_cpu.cpu.genblk3.csr.mcause3_0\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12572_ _05872_ _01003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_184_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13784__A3 _06785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_212_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07999__A1 _02302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11789__S _05336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_200_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14311_ _00165_ net3 mod.u_cpu.rf_ram.memory\[532\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__15337__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11523_ _05144_ mod.u_cpu.rf_ram.memory\[27\]\[0\] _05156_ _05157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_196_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15291_ _00050_ net4 mod.u_scanchain_local.module_data_in\[48\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08660__A2 _02966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_200_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14242_ _00096_ net3 mod.u_cpu.rf_ram.memory\[566\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_183_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14194__B1 _03674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11454_ _05108_ mod.u_cpu.rf_ram.memory\[290\]\[1\] _05103_ _05109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_137_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12744__A1 _05843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_183_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10405_ _04395_ _00313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_11385_ _04377_ _05062_ _05063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_14173_ _07080_ _01396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_152_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14361__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15487__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13124_ _06237_ mod.u_cpu.rf_ram.memory\[359\]\[1\] _06248_ _06251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_139_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10336_ _04347_ _04348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_98_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12413__S _05758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13055_ _06205_ mod.u_cpu.rf_ram.memory\[82\]\[0\] _06206_ _06207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_10267_ _03751_ _04299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__13736__C _06381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_238_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_239_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12006_ _05487_ _05488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_152_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_266_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10198_ _04251_ _03873_ _04252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_254_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07923__B2 _02230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_226_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_207_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_253_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_235_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13957_ _06927_ _06929_ _01331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_46_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08479__A2 _02782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08846__B _02377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_228_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_263_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_250_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12908_ _06086_ mod.u_cpu.rf_ram.memory\[97\]\[1\] _06093_ _06095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_13888_ mod.u_cpu.cpu.immdec.imm30_25\[0\] _06640_ _06877_ _06879_ _06835_ _06880_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_185_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_179_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15627_ _01398_ net3 mod.u_cpu.rf_ram.memory\[8\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2080 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12839_ _05888_ _06048_ _06049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13224__A2 _06326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2091 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_163_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_159_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15558_ _01329_ net3 mod.u_arbiter.i_wb_cpu_dbus_dat\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12283__I0 _05660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08100__A1 _02406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11786__A2 _05335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07534__S0 _01841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14509_ _00363_ net3 mod.u_cpu.rf_ram.memory\[433\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_175_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15489_ _01260_ net3 mod.u_arbiter.i_wb_cpu_dbus_adr\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_163_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08030_ mod.u_cpu.rf_ram.memory\[80\]\[0\] mod.u_cpu.rf_ram.memory\[81\]\[0\] mod.u_cpu.rf_ram.memory\[82\]\[0\]
+ mod.u_cpu.rf_ram.memory\[83\]\[0\] _02249_ _02098_ _02338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__14704__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08403__A2 _02702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_192_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10597__I0 _04523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09981_ _03933_ _04087_ _04097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_254_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14854__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08932_ mod.u_cpu.rf_ram.memory\[535\]\[1\] _03239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__12323__S _05700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13696__C1 _06493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_257_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11010__I1 mod.u_cpu.rf_ram.memory\[360\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_97_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08863_ _02472_ _03169_ _03170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_218_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07914__A1 _02220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07814_ _01719_ _02122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_111_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08794_ _02202_ _03099_ _03100_ _02086_ _03101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_245_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_211_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11849__I0 _05366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10778__S _04645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07745_ _01444_ _02053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_84_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_37_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_226_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07676_ _01962_ mod.u_cpu.rf_ram.memory\[276\]\[0\] _01983_ _01984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09431__I mod.u_cpu.cpu.immdec.imm11_7\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07142__A2 _01440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_213_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07773__S0 _02048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_240_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__14234__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09415_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[28\] _03638_ _03648_ _03649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__09419__A1 _03439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10577__I _04250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_201_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09346_ _03588_ _03590_ _03591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_139_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_194_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12792__I _06017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09277_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[7\] mod.u_cpu.cpu.ctrl.o_ibus_adr\[6\] _03532_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_20_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14384__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08228_ _02534_ _02535_ _02536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_148_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12726__A1 _03885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08159_ _02120_ _02467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11201__I _04879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11170_ _04915_ _00558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_134_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10121_ _04194_ _04195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12329__I1 mod.u_cpu.rf_ram.memory\[184\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_249_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_216_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08158__A1 _02461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10052_ _04146_ _00209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_5634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_88_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4900 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_196_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07905__A1 _02211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_236_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4911 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_236_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4922 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_130_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4933 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14860_ _00714_ net3 mod.u_cpu.rf_ram.memory\[258\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_76_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4944 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_208_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4955 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13829__I1 mod.u_arbiter.i_wb_cpu_rdt\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_180_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4966 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13811_ _06337_ _06811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_235_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4977 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4988 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14791_ _00645_ net3 mod.u_cpu.rf_ram.memory\[292\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_28_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4999 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_169_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08705__I0 mod.u_cpu.rf_ram.memory\[238\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_232_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13742_ _06459_ _06712_ _06747_ _06423_ _06748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__10268__A2 _04133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10954_ _03871_ _04766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_113_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_232_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_204_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08330__A1 _02559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07764__S0 _02070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_189_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13673_ _06683_ _06293_ _06282_ _06294_ _06684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_71_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10885_ _04719_ _04720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_231_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_15412_ _01187_ net3 mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__14727__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12624_ _05907_ mod.u_cpu.rf_ram.memory\[151\]\[1\] _05905_ _05908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XPHY_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__07516__S0 _01823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_200_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11768__A2 _05321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12965__A1 _06135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_200_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15343_ _01118_ net3 mod.u_cpu.rf_ram.memory\[399\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12555_ _05861_ _00997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_185_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_145_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_258_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11506_ _05144_ mod.u_cpu.rf_ram.memory\[282\]\[0\] _05145_ _05146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_184_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15274_ _00032_ net4 mod.u_arbiter.i_wb_cpu_rdt\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__13509__A3 _03260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12486_ _05606_ _05767_ _05817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_172_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14877__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_176_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14225_ _00001_ net3 mod.u_cpu.rf_ram.rdata\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11437_ _04821_ _05089_ _05097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10579__I0 _04506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08397__A1 _02111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13390__A1 _05784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_217_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_193_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14156_ _07067_ _03284_ _07068_ _01391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_11368_ _04766_ _05038_ _05052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_125_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08492__S1 _02666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11940__A2 _05423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13107_ _02284_ _06239_ _06240_ _01170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_140_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10319_ _04311_ _04336_ _04337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_14087_ _07024_ _01366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_11299_ _04978_ mod.u_cpu.rf_ram.memory\[315\]\[0\] _05004_ _05005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_112_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09516__I _03739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09197__I0 mod.u_arbiter.i_wb_cpu_rdt\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_239_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_234_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14190__I0 _07081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_224_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_13038_ _06195_ _01146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_140_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_255_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_187_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10751__I0 _04622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14257__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14989_ _00843_ net3 mod.u_cpu.rf_ram.memory\[29\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_47_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__15502__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_208_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07530_ _01503_ _01838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_19_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08321__A1 _02592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_222_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07461_ _01742_ _01748_ _01767_ _01768_ _01769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_179_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09200_ _03472_ _00028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_210_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07392_ _01497_ _01700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_72_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_188_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12956__A1 _06121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_203_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09131_ _03424_ _03387_ _03427_ _03421_ _00052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_175_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12318__S _05697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08624__A2 _02930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_191_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09062_ _03356_ _03365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_124_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_198_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_147_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10431__A2 _04380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_175_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_200_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_200_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08013_ _01719_ _02321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_116_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13381__A1 _06413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11231__I1 _04954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_235_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09964_ _04085_ _00182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__15032__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09188__I0 mod.u_arbiter.i_wb_cpu_rdt\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10990__I0 _04772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_170_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08915_ _02550_ mod.u_cpu.rf_ram.memory\[526\]\[1\] _03221_ _02515_ _03222_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_09895_ _03829_ _04038_ _04039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09888__A1 _03823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11892__S _05409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_218_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_4229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11695__A1 _04852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08846_ _02365_ _03152_ _02377_ _03153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08560__A1 _01998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_217_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15182__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08777_ _02329_ mod.u_cpu.rf_ram.memory\[118\]\[1\] _03083_ _01916_ _03084_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_2805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_226_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11447__A1 _04831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07728_ _01738_ _01976_ _02035_ _02036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_26_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12495__I0 _05822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09161__I mod.u_arbiter.i_wb_cpu_rdt\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08312__A1 _02592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11998__A2 _05481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_241_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_198_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07659_ _01758_ _01967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_213_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10100__I _03828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10670_ _04568_ _04574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_167_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_159_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__12947__A1 _03500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09329_ _03554_ mod.u_scanchain_local.module_data_in\[52\] _03555_ mod.u_arbiter.i_wb_cpu_dbus_adr\[15\]
+ _03577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_107_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08615__A2 _02921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12340_ _05712_ _00931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_167_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_193_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10973__A3 _03724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12271_ _05665_ _00909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_111_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_209_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_153_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08379__A1 _02561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14010_ _06909_ _06970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_257_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11222_ _04938_ mod.u_cpu.rf_ram.memory\[326\]\[0\] _04949_ _04950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_175_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_218_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_162_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10770__I _04640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11153_ _04896_ mod.u_cpu.rf_ram.memory\[338\]\[1\] _04902_ _04904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_122_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09179__I0 mod.u_arbiter.i_wb_cpu_rdt\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10104_ _04178_ mod.u_cpu.rf_ram.memory\[502\]\[1\] _04181_ _04183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__14172__I0 _07057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11084_ _04857_ _00530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_89_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13675__A2 _06490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15525__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_237_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_14912_ _00766_ net3 mod.u_cpu.rf_ram.memory\[22\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10035_ mod.u_cpu.cpu.immdec.imm11_7\[2\] _03715_ _03717_ _04133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__12722__I1 _05971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_49_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_209_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10733__I0 _04608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_264_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14843_ _00697_ net3 mod.u_cpu.rf_ram.memory\[266\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_124_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_264_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14774_ _00628_ net3 mod.u_cpu.rf_ram.memory\[300\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_189_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11986_ _05474_ _00815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_90_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_205_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_204_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11989__A2 _05475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13725_ _06729_ _06730_ _06731_ _06314_ _06713_ _06732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_95_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10937_ _04753_ mod.u_cpu.rf_ram.memory\[371\]\[0\] _04754_ _04755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_189_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_220_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_232_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_13656_ _06312_ _06392_ _06668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_108_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10868_ _04702_ _04708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_73_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_176_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08843__C _02093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12607_ _04024_ _05896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_157_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_83_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13587_ _03692_ _06614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_223_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10799_ _04660_ _00442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_173_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15326_ _01103_ net3 mod.u_cpu.cpu.state.ibus_cyc vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_118_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_12538_ _02131_ _05849_ _05850_ _00991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_8_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07459__C _01766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_201_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15257_ _00013_ net4 mod.u_arbiter.i_wb_cpu_rdt\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07290__A1 _01561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12469_ _05805_ _00967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__15055__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14208_ _03775_ _07100_ _07101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12166__A2 _05319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15188_ _01041_ net3 mod.u_cpu.rf_ram.memory\[77\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11776__I _05328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14139_ _03980_ _04996_ _07058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_154_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09246__I _03493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07593__A2 _01892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_230_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08700_ _01573_ mod.u_cpu.rf_ram.memory\[198\]\[1\] _03006_ _02212_ _03007_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_09680_ _03875_ _00108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08542__A1 _02091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07345__A2 _01639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08631_ _01818_ _02935_ _02937_ _02938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_95_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_254_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08562_ _01967_ _02868_ _02869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_130_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12477__I0 _05807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_223_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07513_ _01820_ _01821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_120_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13940__B _06914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08493_ mod.u_cpu.rf_ram.memory\[333\]\[1\] _02800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__10101__A1 _04180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_223_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_250_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07444_ _01645_ _01752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_23_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10652__A2 _04437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_241_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10855__I _04640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07375_ _01665_ _01683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_31_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09114_ _03405_ _03413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_149_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09045_ _03253_ _03349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07281__A1 _01446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_191_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_198_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_191_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_209_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13354__A1 _06434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_239_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14422__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15548__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13106__A1 _05948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09156__I mod.u_arbiter.i_wb_cpu_dbus_dat\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09947_ _04073_ mod.u_cpu.rf_ram.memory\[526\]\[0\] _04074_ _04075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__13657__A2 _06668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4004 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_219_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4015 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4026 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09878_ _04023_ mod.u_cpu.rf_ram.memory\[537\]\[0\] _04027_ _04028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__13834__C _03682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14572__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4037 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_213_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4048 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08533__A1 _02225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4059 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08829_ _02411_ _03135_ _03136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_3325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07832__C _02139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12468__I0 _05753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11840_ _03993_ _05371_ _05372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_2624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_227_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1901 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1923 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_214_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_199_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11771_ _03903_ _05325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_1934 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1945 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_207_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_202_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1956 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13510_ _06564_ _06565_ _06566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_214_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10722_ _04608_ mod.u_cpu.rf_ram.memory\[406\]\[1\] _04606_ _04609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_1967 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_214_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14490_ _00344_ net3 mod.u_cpu.rf_ram.memory\[442\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1978 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11840__A1 _03993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1989 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_13441_ _06522_ _01222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__10765__I _04621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_201_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10653_ _04557_ mod.u_cpu.rf_ram.memory\[417\]\[0\] _04562_ _04563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_142_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15078__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08144__S0 _02450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12396__A2 _04335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_220_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13372_ _06292_ _06468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08235__I _01855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10584_ _04233_ _04507_ _04516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_155_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15111_ _00965_ net3 mod.u_cpu.rf_ram.memory\[172\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_177_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07272__A1 _01578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12323_ _05696_ mod.u_cpu.rf_ram.memory\[179\]\[0\] _05700_ _05701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_103_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15042_ _00896_ net3 mod.u_cpu.rf_ram.memory\[197\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_142_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12254_ _05408_ _05650_ _05654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_142_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09013__A2 _03305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_181_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11205_ _04808_ _03986_ _04939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_141_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12185_ _05606_ _05568_ _05607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_123_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_218_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07575__A2 mod.u_cpu.rf_ram.memory\[374\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14915__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14145__I0 _07057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11136_ _04880_ mod.u_cpu.rf_ram.memory\[341\]\[1\] _04891_ _04893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_95_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_231_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11659__A1 _04973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11067_ _04844_ _04845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_110_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xtiny_user_project_120 la_data_out[38] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_62_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08524__A1 _01879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_131 la_data_out[49] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_95_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_142 la_data_out[60] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_5283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_49_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10018_ _03975_ _04118_ _04122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_77_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_236_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xtiny_user_project_153 wbs_dat_o[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_4560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xtiny_user_project_164 wbs_dat_o[14] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_64_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xtiny_user_project_175 wbs_dat_o[25] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__10182__I1 mod.u_cpu.rf_ram.memory\[491\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_149_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14826_ _00680_ net3 mod.u_cpu.rf_ram.memory\[274\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_4593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12220__I _05629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_252_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_205_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14757_ _00611_ net3 mod.u_cpu.rf_ram.memory\[30\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08827__A2 mod.u_cpu.rf_ram.memory\[20\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11969_ _05448_ _05462_ _05463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__11131__I0 _04880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_229_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13820__A2 _06458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_251_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_232_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13708_ _06318_ _06364_ _06713_ _06715_ _06365_ _06716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_44_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_260_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14688_ _00542_ net3 mod.u_cpu.rf_ram.memory\[343\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_220_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13639_ mod.u_cpu.cpu.immdec.imm19_12_20\[0\] _06651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_60_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10675__I _04496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_177_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07160_ _01468_ _01469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_160_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11434__I1 _05065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10398__A1 _02436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14445__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_173_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15309_ _00070_ net4 mod.u_scanchain_local.module_data_in\[66\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_121_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13336__A1 _06423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09177__S _03459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08438__S1 _01995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13887__A2 _06850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_236_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11898__A1 _04973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14595__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10945__I0 _04753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09801_ _03958_ mod.u_cpu.rf_ram.memory\[547\]\[0\] _03970_ _03971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__14136__I0 _07055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_259_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_262_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07993_ _02297_ mod.u_cpu.rf_ram.memory\[108\]\[0\] _02300_ _02301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_141_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09732_ _03915_ _03916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_171_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__12698__I0 _05934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08515__A1 _02759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07949__S0 _02242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_228_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08748__C _01751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09663_ _03763_ _03862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_83_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_255_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08610__S1 _02049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08614_ mod.u_cpu.rf_ram.memory\[148\]\[1\] mod.u_cpu.rf_ram.memory\[149\]\[1\] mod.u_cpu.rf_ram.memory\[150\]\[1\]
+ mod.u_cpu.rf_ram.memory\[151\]\[1\] _02059_ _01723_ _02921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_09594_ _03725_ _03807_ _03808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_70_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_247_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08545_ _01886_ _02852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_42_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08818__A2 mod.u_cpu.rf_ram.memory\[28\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09866__I1 mod.u_cpu.rf_ram.memory\[53\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_251_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10625__A2 _04534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15220__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08476_ mod.u_cpu.rf_ram.memory\[367\]\[1\] _02783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_11_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_211_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_145_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07427_ _01493_ _01724_ _01734_ _01534_ _01735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_17_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_210_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08055__I _01586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07358_ _01665_ _01666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_176_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10389__A1 _04233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09243__A2 _03503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15370__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07289_ mod.u_cpu.rf_ram.memory\[503\]\[0\] _01597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_163_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07894__I _01779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14938__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09028_ _03307_ _03330_ _03251_ _03331_ _03332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_164_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_172_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12925__I1 mod.u_cpu.rf_ram.memory\[379\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08754__A1 _02171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13845__B _06450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_172_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_266_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_172_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13990_ mod.u_arbiter.i_wb_cpu_dbus_dat\[11\] _06954_ _06955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_219_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08506__A1 _02672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12941_ _06117_ _06118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_218_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__13136__I _06252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_219_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_206_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14318__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12872_ _06070_ mod.u_cpu.rf_ram.memory\[409\]\[1\] _06068_ _06071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_234_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14611_ _00465_ net3 mod.u_cpu.rf_ram.memory\[382\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11823_ _05360_ _00766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_61_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15591_ _01362_ net3 mod.u_cpu.rf_ram.memory\[114\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08809__A2 _03088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_233_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13802__A2 _06466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09857__I1 mod.u_cpu.rf_ram.memory\[540\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_214_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_214_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14542_ _00396_ net3 mod.u_cpu.rf_ram.memory\[416\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11754_ _05311_ mod.u_cpu.rf_ram.memory\[238\]\[0\] _05313_ _05314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_183_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_261_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_198_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_261_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08393__C _02606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14468__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_187_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10705_ _04597_ _00411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10495__I _03790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14473_ _00327_ net3 mod.u_cpu.rf_ram.memory\[451\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_14_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11685_ _02273_ _05264_ _05266_ _00722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_186_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_224_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08117__S0 _02391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12369__A2 _04137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13424_ _06510_ _06511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_186_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10636_ _04523_ mod.u_cpu.rf_ram.memory\[420\]\[0\] _04551_ _04552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_167_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13355_ _06450_ _06451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_139_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12416__S _05763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10567_ _01780_ _04503_ _04504_ _00366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_259_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12306_ _05677_ mod.u_cpu.rf_ram.memory\[186\]\[1\] _05687_ _05689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_182_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13286_ _06291_ _06293_ _06384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_170_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10498_ _04459_ _00342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_108_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13869__A2 _06438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15025_ _00879_ net3 mod.u_cpu.rf_ram.memory\[76\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_142_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12916__I1 _05971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12237_ _05642_ _05641_ _05643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_123_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14118__I0 _07043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12541__A2 _05831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12168_ _05322_ _05595_ _05596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_151_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10552__A1 _04360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11119_ _04881_ _00541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07753__B _01632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12099_ _05548_ _00854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_110_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_65_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xtiny_user_project_70 io_out[26] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_232_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5080 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xtiny_user_project_81 io_out[37] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_110_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5091 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_237_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_225_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_92 la_data_out[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_36_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11352__I0 _05032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11990__S _05475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15243__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_266_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_14809_ _00663_ net3 mod.u_cpu.rf_ram.memory\[283\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_18_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_233_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08330_ _02559_ mod.u_cpu.rf_ram.memory\[500\]\[1\] _02636_ _02637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_221_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_205_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08276__A3 _02522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_221_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15393__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08261_ _02533_ mod.u_cpu.rf_ram.memory\[534\]\[0\] _02568_ _02537_ _02569_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_221_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_220_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_123_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07212_ _01519_ _01520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08192_ _02216_ _02500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_193_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07236__A1 _01508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07143_ _01431_ _01423_ _01452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07331__S1 _01638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07647__C _01768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10791__A1 _04242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12125__I _05549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07539__A2 _01846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09784__I0 _03936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12532__A2 _05846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_43_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11591__I0 _05194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__12061__S _05522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07976_ mod.u_cpu.rf_ram.memory\[101\]\[0\] _02284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_56_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09536__I0 _03740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09434__I mod.u_cpu.cpu.immdec.imm11_7\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08478__C _02030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09715_ _03870_ _03883_ _03903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_228_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_216_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11343__I0 _05028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09646_ _03704_ _03819_ _03848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_216_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__14037__A2 _06989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07711__A2 _02011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09577_ _03764_ mod.u_cpu.rf_ram.memory\[571\]\[1\] _03792_ _03794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__13096__I0 _06217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14610__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_215_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13796__A1 _06321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08528_ _01977_ _02817_ _02834_ _02835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_93_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_243_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11271__A2 _04984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08459_ mod.u_cpu.rf_ram.memory\[376\]\[1\] mod.u_cpu.rf_ram.memory\[377\]\[1\] mod.u_cpu.rf_ram.memory\[378\]\[1\]
+ mod.u_cpu.rf_ram.memory\[379\]\[1\] _01957_ _01958_ _02766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_211_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11204__I _04882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_211_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_196_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14760__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_211_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11470_ _05119_ _05120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_168_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_149_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_221_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10421_ _04387_ mod.u_cpu.rf_ram.memory\[455\]\[1\] _04404_ _04406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07227__A1 _01493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_178_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08814__I2 _03119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10082__I0 _04157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13140_ _06260_ _01183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_136_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10352_ _04345_ mod.u_cpu.rf_ram.memory\[466\]\[1\] _04357_ _04359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_87_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_191_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15116__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_183_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13071_ _06216_ _01158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_151_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10283_ _01557_ _04310_ _04312_ _00274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_151_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12022_ _05412_ _05498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_183_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13720__A1 _06726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11874__I _05386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_266_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_266_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__15266__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13973_ _06914_ _06942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_93_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12924_ _06104_ _06105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_111_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12039__A1 _05443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14290__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08750__I1 mod.u_cpu.rf_ram.memory\[105\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_15643_ _01414_ net3 mod.u_cpu.rf_ram.memory\[259\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_62_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12855_ _06058_ _01100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_262_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_222_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11806_ _02237_ _05347_ _05349_ _00760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__13787__A1 _06774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11637__I1 mod.u_cpu.rf_ram.memory\[260\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15574_ _01345_ net3 mod.u_arbiter.i_wb_cpu_dbus_dat\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_61_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12786_ _05998_ mod.u_cpu.rf_ram.memory\[131\]\[1\] _06012_ _06014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_2295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09455__A2 _03681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08889__S1 _02473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14525_ _00379_ net3 mod.u_cpu.rf_ram.memory\[425\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11737_ _05254_ _05301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_203_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_202_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_109_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14456_ _00310_ net3 mod.u_cpu.rf_ram.memory\[45\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11668_ _05253_ _05254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_186_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__14200__A2 _06151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07218__A1 _01517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13407_ _03790_ _06344_ _06500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_174_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10619_ _03773_ _04541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_128_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14387_ _00241_ net3 mod.u_cpu.rf_ram.memory\[494\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11599_ _05199_ mod.u_cpu.rf_ram.memory\[266\]\[0\] _05206_ _05207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_155_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07313__S1 _01570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13338_ _06379_ _06435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08423__I _01914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_192_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_182_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13269_ _06298_ _06367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_131_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08718__A1 _01704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15008_ _00862_ net3 mod.u_cpu.rf_ram.memory\[20\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__13711__A1 _06716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15609__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12514__A2 _05667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11573__I0 _05178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08813__S1 _02267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__11784__I _03917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07830_ _02136_ _02137_ _02138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08298__C _02196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07761_ _02046_ _02068_ _02051_ _02069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_110_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14633__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_256_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09500_ _03725_ _03726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09143__A1 mod.u_arbiter.i_wb_cpu_rdt\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08577__S0 _02020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_225_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10828__A2 _04669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07692_ _01711_ _01999_ _02000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13932__C _03269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09431_ mod.u_cpu.cpu.immdec.imm11_7\[3\] _03662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_266_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_225_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_252_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13778__A1 _06404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13778__B2 _06426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09362_ _03563_ mod.u_scanchain_local.module_data_in\[58\] _03517_ mod.u_arbiter.i_wb_cpu_dbus_adr\[21\]
+ _03604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__14783__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_244_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08313_ mod.u_cpu.rf_ram.memory\[464\]\[1\] mod.u_cpu.rf_ram.memory\[465\]\[1\] mod.u_cpu.rf_ram.memory\[466\]\[1\]
+ mod.u_cpu.rf_ram.memory\[467\]\[1\] _02593_ _02454_ _02620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_178_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09293_ _03528_ _03544_ _03545_ _00050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__12450__A1 _05780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_221_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08244_ mod.u_cpu.rf_ram.memory\[527\]\[0\] _02552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_192_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15139__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_203_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08175_ _02175_ _02483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_165_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08501__S0 _01920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13950__A1 mod.u_arbiter.i_wb_cpu_rdt\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07126_ mod.u_cpu.cpu.decode.op21 _01435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_133_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15289__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_217_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08709__A1 _02594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_153_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08185__A2 _02492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09382__A1 _03564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09164__I _03413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_248_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07959_ _01614_ _02267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_101_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_262_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_216_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09134__A1 _03428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08568__S0 _01957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08001__C _02308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10970_ _04777_ _00496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_21_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_210_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_216_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07696__A1 _01722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08936__C _02518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09629_ _03702_ _03820_ _03835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_244_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_188_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12640_ _05917_ _01026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_70_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07791__S1 _02098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13769__A1 _03670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_188_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12816__I0 _06019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07412__I _01719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_197_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07448__A1 _01728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12571_ _05869_ mod.u_cpu.rf_ram.memory\[15\]\[0\] _05871_ _05872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_141_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_239_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_178_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_197_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14310_ _00164_ net3 mod.u_cpu.rf_ram.memory\[532\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_197_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11522_ _05110_ _03791_ _05156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_156_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07999__A2 mod.u_cpu.rf_ram.memory\[110\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15290_ _00049_ net4 mod.u_scanchain_local.module_data_in\[47\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_184_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_200_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_14241_ _00095_ net3 mod.u_cpu.rf_ram.memory\[567\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11453_ _05107_ _05108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10773__I _03895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14506__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12744__A2 _05986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10404_ _04387_ mod.u_cpu.rf_ram.memory\[458\]\[1\] _04393_ _04395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08243__I _01863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14172_ _07057_ mod.u_cpu.rf_ram.memory\[88\]\[0\] _07079_ _07080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_11384_ _03892_ _04779_ _05062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_164_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10755__A1 _04209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13123_ _01906_ _06248_ _06250_ _01176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_217_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07620__A1 _01925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10335_ _04247_ _04347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_11_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13054_ _03858_ _06193_ _06206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_152_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10266_ _04248_ _04298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_87_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14656__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10507__A1 _04163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12005_ _03773_ _05487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09373__A1 _03489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_266_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10197_ _04250_ _04251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11180__A1 _04379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__11307__I0 _04999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_238_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13956_ mod.u_arbiter.i_wb_cpu_rdt\[2\] _06906_ _06928_ _03438_ _06929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_35_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_207_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_207_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12907_ _06094_ _01116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_13887_ _06823_ _06850_ _06878_ _06423_ _06409_ _06879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_62_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11045__S _04828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_234_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_222_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2070 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09023__B _03268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12838_ _05720_ _06048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_15626_ _01397_ net3 mod.u_cpu.rf_ram.memory\[88\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_185_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2081 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2092 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_250_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12432__A1 _05593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12769_ _06002_ _01070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_15557_ _01328_ net3 mod.u_cpu.rf_ram.memory\[111\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_163_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_203_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_226_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07534__S1 _01763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_175_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10294__I0 _04298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_14508_ _00362_ net3 mod.u_cpu.rf_ram.memory\[433\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_15488_ _01259_ net3 mod.u_arbiter.i_wb_cpu_dbus_adr\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_175_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12035__I1 _05437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14439_ _00293_ net3 mod.u_cpu.rf_ram.memory\[468\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_190_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09249__I _03502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08939__A1 _01464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08153__I _02115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15431__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09987__I0 _04096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13932__A1 _03268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07298__S0 _01605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_183_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13994__I _06910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09980_ _04050_ _04096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_192_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09739__I0 _03890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08931_ _02546_ mod.u_cpu.rf_ram.memory\[532\]\[1\] _03237_ _03238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_88_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13696__B1 _06464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_170_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__15581__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08798__S0 _01561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08862_ mod.u_cpu.rf_ram.memory\[549\]\[1\] _03169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_69_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07914__A2 _02221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07813_ _02110_ _02114_ _02119_ _02120_ _02121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_57_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08793_ _02161_ mod.u_cpu.rf_ram.memory\[76\]\[1\] _03100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_244_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_257_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07744_ _02046_ _02050_ _02051_ _02052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_38_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07678__A1 _01949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_226_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07675_ _01934_ _01982_ _01983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_16_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09414_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[29\] _03648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_52_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07773__S1 _02049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_197_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_164_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_201_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07232__I _01539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09345_ _03542_ _03538_ _03589_ _03585_ _03590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_244_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_205_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10285__I0 _04313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__14529__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09276_ _03528_ _03530_ _03531_ _00047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_138_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08227_ mod.u_cpu.rf_ram.memory\[519\]\[0\] _02535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_193_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_194_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_181_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__12726__A2 _05576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_180_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08158_ _02461_ mod.u_cpu.rf_ram.memory\[550\]\[0\] _02464_ _02465_ _02466_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__14679__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07109_ mod.u_cpu.rf_ram_if.rtrig0 _01418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07602__A1 _01872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08089_ _02302_ mod.u_cpu.rf_ram.memory\[28\]\[0\] _02396_ _02397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_136_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10120_ _03722_ _03726_ _04194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_121_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_255_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10051_ _04140_ mod.u_cpu.rf_ram.memory\[510\]\[1\] _04144_ _04146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_5624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_87_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11162__A1 _04766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4901 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4912 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07905__A2 mod.u_cpu.rf_ram.memory\[210\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_249_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4923 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07756__I2 mod.u_cpu.rf_ram.memory\[138\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_180_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4934 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4945 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_189_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_263_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4956 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14100__A1 _03885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4967 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13810_ _06476_ _06806_ _06809_ _06810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_75_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4978 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14790_ _00644_ net3 mod.u_cpu.rf_ram.memory\[292\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_1_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4989 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_169_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13741_ _06745_ _06746_ _06462_ _06747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_44_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_250_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10953_ _04765_ _00491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_44_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15304__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_186_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_216_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08330__A2 mod.u_cpu.rf_ram.memory\[500\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_204_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07764__S1 _02071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13672_ _06291_ _06683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08238__I _02477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10884_ _04496_ _04719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_232_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_232_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_223_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_15411_ _01186_ net3 mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_71_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12623_ _05873_ _05907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_185_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_197_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08682__B _02988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_157_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08713__S0 _01507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07516__S1 _01821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15342_ _01117_ net3 mod.u_cpu.rf_ram.memory\[97\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_212_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08094__A1 _02348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15454__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12554_ _05855_ mod.u_cpu.rf_ram.memory\[162\]\[0\] _05860_ _05861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_157_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__10976__A1 _04414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11505_ _04868_ _05125_ _05145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_78_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_15273_ _00031_ net4 mod.u_arbiter.i_wb_cpu_rdt\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_32_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_200_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12485_ _05816_ _00972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_7_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14224_ _00000_ net3 mod.u_cpu.rf_ram.rdata\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09969__I0 _04073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11436_ _05045_ _05096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09594__A1 _03725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08397__A2 _02703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14155_ _06057_ _06111_ _07068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10008__I _04090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11367_ _05051_ _00619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_152_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_259_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13106_ _05948_ _06239_ _06240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_3_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10318_ _04172_ _04335_ _04336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_256_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14086_ _06904_ mod.u_cpu.rf_ram.memory\[113\]\[1\] _07022_ _07024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_11298_ _04457_ _04990_ _05004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13319__I _06415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13037_ _06186_ mod.u_cpu.rf_ram.memory\[83\]\[0\] _06194_ _06195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_152_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10249_ _04276_ mod.u_cpu.rf_ram.memory\[481\]\[0\] _04286_ _04287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_266_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_226_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_239_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10751__I1 mod.u_cpu.rf_ram.memory\[401\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07761__B _02051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_187_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14988_ _00842_ net3 mod.u_cpu.rf_ram.memory\[29\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_82_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_240_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_228_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13939_ _06913_ _06914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_208_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08321__A2 _02620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_179_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07460_ _01586_ _01768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_179_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08148__I _02129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_223_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13989__I _06942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_179_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15609_ _01380_ net3 mod.u_cpu.rf_ram.memory\[116\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_50_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07391_ mod.u_cpu.rf_ram.memory\[408\]\[0\] mod.u_cpu.rf_ram.memory\[409\]\[0\] mod.u_cpu.rf_ram.memory\[410\]\[0\]
+ mod.u_cpu.rf_ram.memory\[411\]\[0\] _01697_ _01698_ _01699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_148_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09130_ _03425_ _03426_ _03427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_148_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_202_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09282__B1 _03536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09061_ mod.u_cpu.cpu.csr_imm _03364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__14821__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13205__I0 mod.u_arbiter.i_wb_cpu_rdt\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07832__A1 _02135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_191_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10019__I0 _04117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_191_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08012_ _02283_ _02315_ _02319_ _02308_ _02320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_194_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13905__A1 _06481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08388__A2 mod.u_cpu.rf_ram.memory\[420\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13381__A2 _06461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08632__I0 mod.u_cpu.rf_ram.memory\[184\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_190_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14971__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_170_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09963_ _04073_ mod.u_cpu.rf_ram.memory\[523\]\[0\] _04084_ _04085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_249_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08914_ _02551_ _03220_ _03221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_58_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09894_ _04002_ _04038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_170_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11144__A1 _03809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09888__A2 _04033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_170_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13673__B _06282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08845_ mod.u_cpu.rf_ram.memory\[40\]\[1\] mod.u_cpu.rf_ram.memory\[41\]\[1\] mod.u_cpu.rf_ram.memory\[42\]\[1\]
+ mod.u_cpu.rf_ram.memory\[43\]\[1\] _02349_ _02393_ _03152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12892__A1 _03974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_170_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15327__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08560__A2 mod.u_cpu.rf_ram.memory\[308\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08776_ _01863_ _03082_ _03083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_3529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_261_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07727_ _01977_ _02009_ _02034_ _02035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_150_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_232_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_150_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12644__A1 _05732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08312__A2 _02610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__14351__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_198_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07658_ _01962_ mod.u_cpu.rf_ram.memory\[300\]\[0\] _01965_ _01966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__15477__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_198_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_214_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07589_ mod.u_cpu.rf_ram.memory\[367\]\[0\] _01897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_129_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10258__I0 _04288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09328_ _03574_ _03575_ _03576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_90_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__14149__A1 _03822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09259_ _03517_ _03518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_154_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_126_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09818__S _03981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12270_ _05660_ mod.u_cpu.rf_ram.memory\[192\]\[1\] _05663_ _05665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_138_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_181_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11221_ _04812_ _04945_ _04949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_49_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08379__A2 _02682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_218_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_150_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_253_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09040__A3 _03259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11152_ _04903_ _00552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_161_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09179__I1 mod.u_arbiter.i_wb_cpu_dbus_dat\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_175_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10103_ _04182_ _00224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_1_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11083_ _04843_ mod.u_cpu.rf_ram.memory\[34\]\[0\] _04856_ _04857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_5421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_191_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14911_ _00765_ net3 mod.u_cpu.rf_ram.memory\[230\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10034_ _03662_ _03665_ _03753_ _04132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XTAP_5454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12978__I _03268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_208_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10733__I1 mod.u_cpu.rf_ram.memory\[404\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08551__A2 mod.u_cpu.rf_ram.memory\[316\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14842_ _00696_ net3 mod.u_cpu.rf_ram.memory\[266\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_4753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_217_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11985_ _05464_ mod.u_cpu.rf_ram.memory\[216\]\[1\] _05472_ _05474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_14773_ _00627_ net3 mod.u_cpu.rf_ram.memory\[301\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_251_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_232_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10497__I0 _04453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13724_ _06382_ _06493_ _06731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_90_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10936_ _04352_ _04733_ _04754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_90_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10110__A2 _04185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_231_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_205_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14844__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13655_ _06304_ _06666_ _06667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_32_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12419__S _05763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10867_ _04707_ _00463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_220_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08067__A1 _02356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12606_ _05895_ _01014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13060__A1 _05948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_31_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13586_ _06613_ _01276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_34_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_12_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10798_ mod.u_cpu.rf_ram.memory\[393\]\[0\] _04658_ _04659_ _04660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XPHY_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12537_ _05642_ _05849_ _05850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_15325_ mod.u_cpu.cpu.o_wdata0 net3 mod.u_cpu.rf_ram_if.wdata0_r vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_173_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14994__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_15256_ _00012_ net4 mod.u_arbiter.i_wb_cpu_rdt\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12468_ _05753_ mod.u_cpu.rf_ram.memory\[419\]\[0\] _05804_ _05805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_138_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11419_ _04539_ _05020_ _05085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_14207_ _03895_ _05210_ _07100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_193_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15187_ _01040_ net3 mod.u_cpu.rf_ram.memory\[142\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_125_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12399_ _05745_ mod.u_cpu.rf_ram.memory\[479\]\[1\] _05750_ _05752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_119_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11374__A1 _05022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09031__A3 _01452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09527__I _03750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10421__I0 _04387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14138_ _06577_ _07057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_98_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14224__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13115__A2 _03986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14069_ mod.u_arbiter.i_wb_cpu_rdt\[31\] _06940_ _07013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_140_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input4_I io_in[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_228_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_255_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_227_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08542__A2 _02848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08630_ _02097_ _02936_ _02937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__14374__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_243_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08561_ mod.u_cpu.rf_ram.memory\[311\]\[1\] _02868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_130_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_214_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__12626__A1 _05494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_208_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13823__B1 _06812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07512_ _01523_ _01820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_223_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08492_ mod.u_cpu.rf_ram.memory\[328\]\[1\] mod.u_cpu.rf_ram.memory\[329\]\[1\] mod.u_cpu.rf_ram.memory\[330\]\[1\]
+ mod.u_cpu.rf_ram.memory\[331\]\[1\] _01920_ _02666_ _02799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_165_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07443_ _01750_ _01751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_165_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_210_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_211_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11233__S _04956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_206_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07374_ _01681_ _01682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07510__I _01657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09113_ mod.u_arbiter.i_wb_cpu_ack _03412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_109_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12128__I _05422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_175_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07805__A1 _01673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_198_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10660__I0 _04560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09044_ _03257_ _03296_ _03319_ _03347_ _03348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_159_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09558__A1 _03700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_190_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13106__A2 _06239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09946_ _03886_ _04062_ _04074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_89_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14717__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_225_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4005 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4016 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07416__S0 _01722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12865__A1 _06063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4027 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09877_ _03996_ _04026_ _04027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4038 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_4049 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08384__I2 mod.u_cpu.rf_ram.memory\[418\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08828_ mod.u_cpu.rf_ram.memory\[23\]\[1\] _03135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_161_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_248_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_173_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08759_ _02352_ _03062_ _03065_ _02361_ _03066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_2614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_233_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__14867__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09089__A3 _03389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1902 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10479__I0 _04430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1913 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_260_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11770_ _05324_ _00749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08297__A1 _02191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_199_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_198_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1924 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_207_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_214_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_213_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_199_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1946 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_199_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10721_ _04578_ _04608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1957 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1968 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12239__S _05641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11840__A2 _05371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1979 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_186_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13440_ _03520_ _06519_ _06520_ _03524_ _06522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_139_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10652_ _04285_ _04437_ _04562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_13_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07420__I _01604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_181_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08144__S1 _02451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09797__A1 _03788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_221_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_13371_ _06463_ _06448_ _06465_ _06466_ _06467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_139_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10583_ _04515_ _00371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_210_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15110_ _00964_ net3 mod.u_cpu.rf_ram.memory\[172\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12322_ _05037_ _05686_ _05700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_127_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14247__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_181_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15041_ _00895_ net3 mod.u_cpu.rf_ram.memory\[119\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12253_ _05653_ _00903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_182_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11204_ _04882_ _04938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_141_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08251__I _01757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_190_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_12184_ _03909_ _05606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_134_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_214_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11135_ _04892_ _00546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__14397__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11108__A1 _04873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12156__I0 _05583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15642__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_237_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11066_ _03990_ _04844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_77_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xtiny_user_project_110 la_data_out[28] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__11659__A2 _05120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_209_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xtiny_user_project_121 la_data_out[39] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_132 la_data_out[50] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_264_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08524__A2 mod.u_cpu.rf_ram.memory\[342\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10017_ _04121_ _00199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_5284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xtiny_user_project_143 la_data_out[61] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_76_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_237_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xtiny_user_project_154 wbs_dat_o[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_114_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xtiny_user_project_165 wbs_dat_o[15] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_4561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09082__I net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_209_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_176 wbs_dat_o[26] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_149_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14825_ _00679_ net3 mod.u_cpu.rf_ram.memory\[275\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_4583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12608__A1 _05896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_184_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13805__B1 _06779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11117__I _04879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14756_ _00610_ net3 mod.u_cpu.rf_ram.memory\[30\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3893 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11968_ _04025_ _05433_ _05462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_91_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11131__I1 mod.u_cpu.rf_ram.memory\[342\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08854__C _01695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13707_ _06683_ _06667_ _06714_ _06493_ _06406_ _06715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_189_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10919_ _04728_ mod.u_cpu.rf_ram.memory\[374\]\[0\] _04742_ _04743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_60_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13408__I0 _06351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11899_ _05413_ mod.u_cpu.rf_ram.memory\[225\]\[0\] _05414_ _05415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_225_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_14687_ _00541_ net3 mod.u_cpu.rf_ram.memory\[344\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_220_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15022__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13638_ _06641_ _06648_ _06650_ _01291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07330__I _01637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08835__I0 mod.u_cpu.rf_ram.memory\[52\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13569_ _03692_ _06604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_118_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_199_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10398__A2 _04390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15308_ _00069_ net4 mod.u_scanchain_local.module_data_in\[65\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_118_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08460__A1 _01956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_173_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15172__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13336__A2 _06430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15239_ _01092_ net3 mod.u_cpu.rf_ram.memory\[124\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_99_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09257__I _03495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08161__I _02143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09800_ _03948_ _03969_ _03970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_99_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07992_ _02298_ _02299_ _02300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_101_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09731_ _03738_ _03915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07933__C _02168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_189_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12847__A1 _02080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13895__I0 _06581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08515__A2 _02818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07949__S1 _02172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09662_ _03861_ _00104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_228_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08613_ _02053_ _02919_ _02920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_209_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09593_ _03718_ _03806_ _03807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_215_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_209_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13647__I0 mod.u_arbiter.i_wb_cpu_rdt\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11027__I _03898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08544_ _02295_ _02847_ _02850_ _01492_ _02851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_242_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_224_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_247_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_208_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08475_ _02022_ mod.u_cpu.rf_ram.memory\[364\]\[1\] _02781_ _02782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_211_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12059__S _05522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_165_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07426_ _01703_ _01727_ _01733_ _01529_ _01734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_196_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_206_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_149_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15515__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07357_ _01499_ _01665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_137_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_191_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07288_ _01556_ mod.u_cpu.rf_ram.memory\[500\]\[0\] _01595_ _01596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_108_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09027_ _03254_ _03331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_191_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10307__S _04328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_191_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_254_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_191_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12386__I0 _05731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08203__A1 _02509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07637__S0 _01774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_176_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09951__A1 _01463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_266_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_219_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_172_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09929_ _04061_ _00171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12689__I1 _05950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08506__A2 _02812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09703__A1 _03724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_246_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_213_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12940_ mod.u_arbiter.i_wb_cpu_rdt\[14\] mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat\[14\]
+ _06116_ _06117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_3101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_219_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12871_ _06018_ _06070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_2422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15045__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14610_ _00464_ net3 mod.u_cpu.rf_ram.memory\[382\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11822_ _05342_ mod.u_cpu.rf_ram.memory\[22\]\[0\] _05359_ _05360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_3189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_261_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15590_ _01361_ net3 mod.u_cpu.rf_ram.memory\[114\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_60_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_199_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_199_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11753_ _05312_ _05301_ _05313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_60_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_14541_ _00395_ net3 mod.u_cpu.rf_ram.memory\[417\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_202_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_187_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10704_ _04593_ mod.u_cpu.rf_ram.memory\[40\]\[1\] _04595_ _04597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_42_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11684_ _05265_ _05264_ _05266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08690__A1 _02578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14472_ _00326_ net3 mod.u_cpu.rf_ram.memory\[451\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_201_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_174_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08117__S1 _01552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15195__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10635_ _04272_ _04534_ _04551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_13423_ _06509_ _06510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_167_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13354_ _06434_ _06435_ _06450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_182_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10566_ _04439_ _04503_ _04504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_155_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12305_ _05688_ _00920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_182_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13285_ _06367_ _06382_ _06383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_142_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11329__A1 _04741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10497_ _04453_ mod.u_cpu.rf_ram.memory\[443\]\[0\] _04458_ _04459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12377__I0 _05729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15024_ _00878_ net3 mod.u_cpu.rf_ram.memory\[76\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_170_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12236_ _03944_ _05642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_5_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12167_ _05593_ _05594_ _05595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_123_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__13755__C _06759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11118_ _04880_ mod.u_cpu.rf_ram.memory\[344\]\[1\] _04877_ _04881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_116_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_231_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12098_ _05539_ mod.u_cpu.rf_ram.memory\[67\]\[0\] _05547_ _05548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_1_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xtiny_user_project_60 io_out[16] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_7_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5070 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11049_ _04827_ mod.u_cpu.rf_ram.memory\[354\]\[0\] _04832_ _04833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xtiny_user_project_71 io_out[27] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_65_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_82 la_data_out[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_265_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5081 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xtiny_user_project_93 la_data_out[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_5092 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07325__I _01494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_266_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_4380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07800__S0 _02106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_237_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_252_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14808_ _00662_ net3 mod.u_cpu.rf_ram.memory\[283\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_224_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_52_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_229_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09540__I _03762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08584__C _02005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_205_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14412__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14739_ _00593_ net3 mod.u_cpu.rf_ram.memory\[318\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__15538__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_178_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_205_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08260_ _02566_ _02567_ _02568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08681__A1 _02632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07211_ _01518_ _01519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08191_ _02456_ mod.u_cpu.rf_ram.memory\[572\]\[0\] _02498_ _02499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_119_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07995__I _01862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07142_ _01432_ _01440_ _01451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_9_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__14562__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10615__I0 _04537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_203_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07236__A2 mod.u_cpu.rf_ram.memory\[460\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08433__A1 _02654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_236_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_160_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_259_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_173_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_248_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11591__I1 mod.u_cpu.rf_ram.memory\[268\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08759__C _02361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07975_ _02212_ _02283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_75_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_228_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09536__I1 mod.u_cpu.rf_ram.memory\[574\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09714_ _03766_ _03902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__15068__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_210_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11343__I1 mod.u_cpu.rf_ram.memory\[308\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_255_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09645_ _03739_ _03847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_132_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07172__A1 mod.u_cpu.cpu.immdec.imm24_20\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09576_ _03793_ _00086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_167_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_243_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08527_ _02822_ _02824_ _02040_ _02833_ _02834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14068__I _03309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_196_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_212_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_208_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_212_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08458_ _02759_ _02760_ _02763_ _02764_ _02765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__14905__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_180_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_51_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_212_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07409_ _01716_ _01717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_149_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08389_ mod.u_cpu.rf_ram.memory\[423\]\[1\] _02696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__11559__A1 _05047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_221_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13700__I _06655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10420_ _01521_ _04404_ _04405_ _00318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__07227__A2 _01502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08424__A1 _02611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08814__I3 _03120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10351_ _04358_ _00296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_100_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09826__S _03987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13070_ _06205_ mod.u_cpu.rf_ram.memory\[81\]\[0\] _06215_ _06216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_124_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10282_ _04311_ _04310_ _04312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_105_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12021_ _05497_ _00827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_133_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_219_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13720__A2 _06314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11731__A1 _05047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_183_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07786__I0 mod.u_cpu.rf_ram.memory\[184\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_250_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08669__C _01723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_266_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_247_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13972_ _03446_ _06911_ _06919_ _05798_ _06941_ _01334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_59_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07538__I0 _01839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14435__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_12923_ _06017_ _06104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_185_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_234_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_207_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13083__S _06224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_206_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15642_ _01413_ net3 mod.u_cpu.rf_ram.memory\[269\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12854_ _06057_ mod.u_cpu.rf_ram_if.rreq_r _06058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_146_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_222_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11098__I0 _04862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11805_ _05348_ _05347_ _05349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_2274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15573_ _01344_ net3 mod.u_arbiter.i_wb_cpu_dbus_dat\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_215_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12785_ _06013_ _01075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_226_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11798__A1 _05343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_261_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_187_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14524_ _00378_ net3 mod.u_cpu.rf_ram.memory\[425\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__14585__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08663__A1 _02711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11736_ _03871_ _05300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_202_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_203_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_230_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10470__A1 _04439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14455_ _00309_ net3 mod.u_cpu.rf_ram.memory\[460\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11667_ _04226_ _05252_ _05253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_30_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_161_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13406_ _04223_ _06358_ _06498_ _06499_ _01210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_128_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07218__A2 mod.u_cpu.rf_ram.memory\[454\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08415__A1 _01459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10618_ _04539_ _04447_ _04540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11598_ _04792_ _05191_ _05206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_190_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14386_ _00240_ net3 mod.u_cpu.rf_ram.memory\[494\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_183_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_259_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12226__I _05634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13337_ _06125_ _06434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_10549_ _04492_ _00360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_115_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_196_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11970__A1 _02203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13268_ _06318_ _06364_ _06365_ _06366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_143_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_237_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_15007_ _00861_ net3 mod.u_cpu.rf_ram.memory\[210\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08718__A2 _03024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11022__I0 _04803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12219_ _03726_ _04226_ _05629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_68_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13199_ _06305_ _06306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__15210__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09391__A2 _03615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07760_ mod.u_cpu.rf_ram.memory\[152\]\[0\] mod.u_cpu.rf_ram.memory\[153\]\[0\] mod.u_cpu.rf_ram.memory\[154\]\[0\]
+ mod.u_cpu.rf_ram.memory\[155\]\[0\] _02066_ _02067_ _02068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_96_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_237_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09143__A2 _03436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08577__S1 _01995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07691_ mod.u_cpu.rf_ram.memory\[285\]\[0\] _01999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__15360__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_253_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11506__S _05145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09430_ _03659_ _03402_ _03493_ _03660_ _03661_ _00073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_24_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10410__S _04397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_225_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14928__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11089__I0 _04843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09361_ _03602_ _03599_ _03603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__13778__A2 _06744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_206_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08312_ _02592_ _02610_ _02618_ _01678_ _02619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_177_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08654__A1 _02110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09292_ _03535_ mod.u_scanchain_local.module_data_in\[47\] _03536_ mod.u_arbiter.i_wb_cpu_dbus_adr\[10\]
+ _03545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_220_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_178_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08243_ _01863_ _02551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_177_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12589__I0 _05869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08174_ _02478_ mod.u_cpu.rf_ram.memory\[556\]\[0\] _02481_ _02482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_174_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07125_ mod.u_cpu.cpu.genblk3.csr.o_new_irq _01434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_192_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08501__S1 _02666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14308__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09206__I0 mod.u_arbiter.i_wb_cpu_rdt\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08709__A2 _03012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11713__A1 _05283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_251_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08489__C _02677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09382__A2 _03617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_251_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14458__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_229_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_214_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_210_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07958_ _02058_ _02266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_169_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09134__A2 _03387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_229_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08568__S1 _01958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07889_ _01519_ _02197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_216_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_216_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09628_ _03766_ _03834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_56_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_249_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_216_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_71_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09559_ _03778_ _03779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_102_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_231_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_231_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11215__I _04905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_168_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12570_ _05870_ _04913_ _05871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_212_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08645__A1 _02110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07448__A2 mod.u_cpu.rf_ram.memory\[420\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_196_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11521_ _05155_ _00669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_212_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_196_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_211_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_200_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11151__S _04902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11452_ _05106_ _05107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_183_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14240_ _00094_ net3 mod.u_cpu.rf_ram.memory\[567\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_149_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14194__A2 _03389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10204__A1 _04255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10403_ _04394_ _00312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_14171_ _03804_ _05397_ _07079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11383_ _05061_ _00625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_178_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_256_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15233__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10755__A2 _04623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13122_ _06249_ _06248_ _06250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_124_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10334_ _04346_ _00291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_124_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07620__A2 mod.u_cpu.rf_ram.memory\[318\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_180_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11885__I _05105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13053_ _06204_ _06205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_180_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10265_ _04297_ _00271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_79_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12004_ _03834_ _04984_ _05486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_152_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_191_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10196_ _03808_ _04250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_39_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07384__A1 _01678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15383__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11180__A2 _04779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_266_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_219_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12504__I0 _05827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09125__A2 _03415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_235_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13955_ _06910_ _06928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_47_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_235_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_185_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07526__I3 _01831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12906_ _06088_ mod.u_cpu.rf_ram.memory\[97\]\[0\] _06093_ _06094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__13209__A1 _06117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_207_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13886_ _06382_ _06285_ _06871_ _06441_ _06878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__09090__I _03390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_262_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_207_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2060 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15625_ _01396_ net3 mod.u_cpu.rf_ram.memory\[88\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_146_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12837_ _06047_ _05788_ _01093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_2071 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2082 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2093 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10818__I0 _04663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15556_ _01327_ net3 mod.u_cpu.rf_ram.memory\[111\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08636__A1 _01836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12432__A2 _05438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12768_ _05998_ mod.u_cpu.rf_ram.memory\[134\]\[1\] _06000_ _06002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_202_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_230_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14507_ _00361_ net3 mod.u_cpu.rf_ram.memory\[434\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11719_ _05221_ _05289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_159_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15487_ _01258_ net3 mod.u_arbiter.i_wb_cpu_dbus_adr\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_187_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12699_ _05957_ _01045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_238_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_14438_ _00292_ net3 mod.u_cpu.rf_ram.memory\[468\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07478__C _01785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08939__A2 _01465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13932__A2 mod.u_cpu.cpu.bufreg.lsb\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09987__I1 mod.u_cpu.rf_ram.memory\[51\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14369_ _00223_ net3 mod.u_cpu.rf_ram.memory\[503\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07298__S1 _01570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11794__I1 _05230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_196_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_157_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14600__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_192_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08930_ _02509_ _03236_ _03237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_115_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13696__B2 _06682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08798__S1 _01714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08861_ mod.u_cpu.rf_ram.memory\[544\]\[1\] mod.u_cpu.rf_ram.memory\[545\]\[1\] mod.u_cpu.rf_ram.memory\[546\]\[1\]
+ mod.u_cpu.rf_ram.memory\[547\]\[1\] _02450_ _02451_ _03168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_96_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_258_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_233_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07812_ _01716_ _02120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_96_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08792_ mod.u_cpu.rf_ram.memory\[77\]\[1\] _03099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_123_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13448__A1 mod.u_cpu.cpu.ctrl.o_ibus_adr\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14750__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07743_ _01661_ _02051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_211_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07674_ mod.u_cpu.rf_ram.memory\[277\]\[0\] _01982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_38_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_203_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07678__A2 _01985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07513__I _01820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15106__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09413_ _03623_ _03646_ _03647_ _00070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_252_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_198_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09344_ _03570_ _03559_ _03589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__13620__A1 _05164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_178_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_240_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_221_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10434__A1 _01512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11482__I0 _05128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_178_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09275_ _03516_ mod.u_scanchain_local.module_data_in\[44\] _03518_ mod.u_arbiter.i_wb_cpu_dbus_adr\[7\]
+ _03531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_32_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_148_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08226_ _02216_ _02534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__15256__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_194_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08157_ _01747_ _02465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_193_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13923__A2 _06899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09978__I1 _03929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08088_ _02369_ _02395_ _02396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07602__A2 _01902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14280__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10315__S _04332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13687__A1 _06292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10050_ _04145_ _00208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_121_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08012__C _02308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11162__A2 _04906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_248_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4902 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_102_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4913 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4924 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_236_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4935 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4946 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_180_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09107__A2 _03406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4957 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_217_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__14100__A2 _07014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4968 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4979 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_217_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_90_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13740_ _06470_ _06425_ _06458_ _06746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_113_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08866__A1 _02462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10952_ _04756_ mod.u_cpu.rf_ram.memory\[36\]\[1\] _04763_ _04765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_244_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_251_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_13671_ _06670_ _06682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_147_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10883_ _04718_ _00468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_204_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_15410_ _01185_ net3 mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_262_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_189_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_12622_ _05906_ _01019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08618__A1 _01849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08682__C _01638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_15341_ _01116_ net3 mod.u_cpu.rf_ram.memory\[97\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08713__S1 _01763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_197_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12553_ _05408_ _05757_ _05860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_185_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08094__A2 _02394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_200_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11504_ _05143_ _05144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_157_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_200_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15272_ _00029_ net4 mod.u_arbiter.i_wb_cpu_rdt\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_71_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__14167__A2 _07075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_185_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12484_ _05807_ mod.u_cpu.rf_ram.memory\[449\]\[1\] _05814_ _05816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_138_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14223_ _00079_ net3 mod.u_cpu.rf_ram.memory\[9\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_172_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14623__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11435_ _05095_ _00643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13914__A2 _06892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09043__A1 _03325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12705__S _05959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11366_ _05050_ mod.u_cpu.rf_ram.memory\[305\]\[1\] _05048_ _05051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09594__A2 _03807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14154_ _06063_ _07067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_98_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13105_ _04107_ _05640_ _06239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_10317_ _04308_ _04335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_152_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11297_ _05003_ _00597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13678__A1 _06421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14085_ _07023_ _01365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__14773__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09085__I _03385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09346__A2 _03590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10248_ _04285_ _04137_ _04286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_13036_ _05732_ _06193_ _06194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_26_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_234_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__13536__S _06584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10179_ _04237_ _00245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_66_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12440__S _05777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_266_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08857__C _01739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15129__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14987_ _00841_ net3 mod.u_cpu.rf_ram.memory\[62\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_93_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13335__I _06431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13150__I0 mod.u_arbiter.i_wb_cpu_rdt\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08857__A1 _02102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13938_ _05800_ _06909_ _06913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_35_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13850__A1 _06472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_235_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_263_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_234_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_223_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13869_ _06694_ _06438_ _06664_ _06283_ _06862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_23_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15608_ _01379_ net3 mod.u_cpu.rf_ram.memory\[116\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__15279__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_250_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08609__A1 _02040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07390_ _01500_ _01698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_195_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_222_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_203_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11464__I0 _05114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15539_ _01310_ net3 mod.u_cpu.cpu.immdec.imm24_20\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__14166__I _06046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_203_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09282__A1 _03535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09060_ _01429_ _03363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_176_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08164__I _02329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08011_ _02316_ mod.u_cpu.rf_ram.memory\[126\]\[0\] _02318_ _02306_ _02319_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_129_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13905__A2 _06660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12615__S _05901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_190_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_200_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07596__A1 _01759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09962_ _03911_ _04062_ _04084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12716__I0 _05963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08913_ mod.u_cpu.rf_ram.memory\[527\]\[1\] _03220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09893_ _04037_ _00159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07348__A1 _01483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11144__A2 _03980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08844_ _02578_ _03147_ _03150_ _02660_ _03151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_97_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12892__A2 _06048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_257_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10869__I _04708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08775_ mod.u_cpu.rf_ram.memory\[119\]\[1\] _03082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_38_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__13141__I0 mod.u_arbiter.i_wb_cpu_rdt\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_175_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_254_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07726_ _01740_ _02019_ _02033_ _02034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_84_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07243__I _01550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09896__I0 _04023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13841__A1 _05787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_226_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_214_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_214_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_214_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_198_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_253_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07657_ _01963_ _01964_ _01965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_26_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_207_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_214_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_198_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07588_ _01893_ mod.u_cpu.rf_ram.memory\[364\]\[0\] _01895_ _01896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_142_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10407__A1 _03714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_179_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14646__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09327_ _03569_ _03560_ _03575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_179_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14149__A2 _05254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09258_ _03407_ _03517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_182_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08209_ _02476_ _02512_ _02516_ _02489_ _02517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_138_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09189_ _03466_ _00023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09025__A1 _01428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08459__S0 _01957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14796__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11220_ _04948_ _00575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_257_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07587__A1 _01759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09040__A4 _03343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11151_ _04901_ mod.u_cpu.rf_ram.memory\[338\]\[0\] _04902_ _04903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_122_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09119__B _03417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10102_ _04162_ mod.u_cpu.rf_ram.memory\[502\]\[0\] _04181_ _04182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_150_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11082_ _04808_ _03975_ _04856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_27_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14910_ _00764_ net3 mod.u_cpu.rf_ram.memory\[230\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_153_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10033_ _04131_ _00205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_5444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_249_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_216_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_4721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_49_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_5466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08677__C _02597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_263_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14841_ _00695_ net3 mod.u_cpu.rf_ram.memory\[267\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_75_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_5499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13132__I0 mod.u_arbiter.i_wb_cpu_rdt\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14772_ _00626_ net3 mod.u_cpu.rf_ram.memory\[301\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_91_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11984_ _05473_ _00814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__15421__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13832__A1 _05790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07153__I _01461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_245_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_217_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_216_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13723_ _06362_ _06668_ _06293_ _06730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10646__A1 _04281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10935_ _04694_ _04753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_264_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_147_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_232_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13654_ _06298_ _06299_ _06666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_140_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_220_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10866_ _04698_ mod.u_cpu.rf_ram.memory\[383\]\[1\] _04705_ _04707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_204_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_34_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_12605_ _05891_ mod.u_cpu.rf_ram.memory\[154\]\[1\] _05893_ _05895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__15571__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13585_ mod.u_arbiter.i_wb_cpu_dbus_adr\[25\] mod.u_arbiter.i_wb_cpu_dbus_adr\[26\]
+ _06609_ _06613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_197_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13060__A2 _06209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10797_ _04527_ _04644_ _04659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_185_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__10949__A2 _03961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11071__A1 _04845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_15324_ _01102_ net3 mod.u_cpu.rf_ram_if.rdata1 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_157_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12536_ _05226_ _05438_ _05849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_185_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_200_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15255_ _00011_ net4 mod.u_arbiter.i_wb_cpu_rdt\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09016__A1 mod.u_cpu.cpu.state.o_cnt_r\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12435__S _05774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12467_ _05649_ _04437_ _05804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13899__A1 _01453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14206_ _06047_ _07073_ _01411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_11418_ _05084_ _00637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_125_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15186_ _01039_ net3 mod.u_cpu.rf_ram.memory\[142\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_158_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12398_ _01562_ _05750_ _05751_ _00950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__11374__A2 _05055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_153_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_193_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14137_ _07056_ _01384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_11349_ _05037_ _05038_ _05039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_153_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08870__S0 _02472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13774__B _06643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14068_ _03309_ _07012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_234_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13019_ _06107_ mod.u_cpu.rf_ram.memory\[10\]\[0\] _06182_ _06183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12170__S _05595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14519__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_239_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_55_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07491__C _01785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_236_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08560_ _01998_ mod.u_cpu.rf_ram.memory\[308\]\[1\] _02866_ _02867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08159__I _02120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09878__I0 _04023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_208_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_223_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07511_ _01506_ _01819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08491_ _01848_ _02777_ _02797_ _02798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__14669__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_235_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07502__A1 _01807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07998__I _01569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07442_ _01749_ _01750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_251_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_167_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_245_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07373_ _01509_ _01681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_195_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11313__I _04951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09112_ _03404_ _03408_ _03411_ _00019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_164_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13949__B _06919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_191_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09043_ _03325_ _03326_ _01394_ _03332_ _03346_ _03347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_163_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14000__A1 mod.u_arbiter.i_wb_cpu_dbus_dat\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07666__C _01812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07569__A1 _01759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08230__A2 mod.u_cpu.rf_ram.memory\[518\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08081__I2 mod.u_cpu.rf_ram.memory\[14\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08861__S0 _02450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09945_ _04050_ _04073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_132_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_213_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08778__B _03084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09876_ _04025_ _04026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_4006 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07416__S1 _01723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10176__I0 _04217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4017 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12865__A2 _06065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15444__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4028 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_245_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_219_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4039 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08827_ _02316_ mod.u_cpu.rf_ram.memory\[20\]\[1\] _03133_ _03134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_3305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10876__A1 _04307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_261_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08069__I _01551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08758_ _02204_ mod.u_cpu.rf_ram.memory\[102\]\[1\] _03064_ _02359_ _03065_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_2615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13814__A1 _06810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09869__I0 _04001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_241_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_227_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09089__A4 mod.u_cpu.cpu.state.o_cnt_r\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11676__I0 _05243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_214_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07709_ _01722_ mod.u_cpu.rf_ram.memory\[262\]\[0\] _02016_ _01970_ _02017_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__10479__I1 mod.u_cpu.rf_ram.memory\[446\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1903 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1914 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08297__A2 mod.u_cpu.rf_ram.memory\[454\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15594__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08689_ _02202_ _02994_ _02995_ _02093_ _02996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_53_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1925 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1936 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_199_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10720_ _04607_ _00416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1947 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_214_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1958 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1969 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_246_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10651_ _04561_ _00393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_167_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_210_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11053__A1 _04285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13370_ _06369_ _06466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_166_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09797__A2 _03966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10582_ _04514_ mod.u_cpu.rf_ram.memory\[42\]\[1\] _04512_ _04515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_103_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12321_ _05699_ _00925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_214_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_142_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_194_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09628__I _03766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15040_ _00894_ net3 mod.u_cpu.rf_ram.memory\[119\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_177_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12252_ _05635_ mod.u_cpu.rf_ram.memory\[195\]\[1\] _05651_ _05653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_154_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_218_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12553__A1 _05408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11203_ _04937_ _00569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_12183_ _05604_ _05605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_163_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11134_ _04883_ mod.u_cpu.rf_ram.memory\[341\]\[0\] _04891_ _04892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_1_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07980__A1 _02136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11065_ _04802_ _04843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_77_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xtiny_user_project_100 la_data_out[18] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_237_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_111 la_data_out[29] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_5263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xtiny_user_project_122 la_data_out[40] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_95_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10016_ _04115_ mod.u_cpu.rf_ram.memory\[515\]\[1\] _04119_ _04121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_5274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xtiny_user_project_133 la_data_out[51] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_4540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_114_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_49_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_144 la_data_out[62] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_97_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14811__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xtiny_user_project_155 wbs_dat_o[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_76_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_237_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xtiny_user_project_166 wbs_dat_o[16] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_64_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_177 wbs_dat_o[27] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_218_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14824_ _00678_ net3 mod.u_cpu.rf_ram.memory\[275\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_4573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_4584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13805__A1 _06468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12608__A2 _05882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_264_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_251_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_151_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14755_ _00609_ net3 mod.u_cpu.rf_ram.memory\[310\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3894 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11967_ _05461_ _00809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_45_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13706_ _06669_ _06714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_264_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_220_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_205_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10918_ _04741_ _04733_ _04742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_233_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__14961__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14686_ _00540_ net3 mod.u_cpu.rf_ram.memory\[344\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_32_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11898_ _04973_ _05401_ _05414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07611__I _01743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_220_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_149_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13637_ mod.u_cpu.cpu.immdec.imm31 _06649_ _06650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_158_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10849_ _04693_ _00459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_201_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_125_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13568_ _06603_ _01268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08835__I1 mod.u_cpu.rf_ram.memory\[53\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15307_ _00068_ net4 mod.u_scanchain_local.module_data_in\[64\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__15317__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_199_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12519_ _05838_ _00984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_200_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_173_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08460__A2 _02766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13499_ _06539_ _06558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_117_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09538__I _03732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_246_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15238_ _01091_ net3 mod.u_cpu.rf_ram.memory\[124\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_173_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13592__I0 mod.u_arbiter.i_wb_cpu_dbus_adr\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15169_ _01022_ net3 mod.u_cpu.rf_ram.memory\[150\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__14341__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__15467__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07991_ mod.u_cpu.rf_ram.memory\[109\]\[0\] _02299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_80_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11509__S _05145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07971__A1 _01739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09730_ _03914_ _00119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10158__I0 _04215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_228_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_227_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09661_ _03847_ mod.u_cpu.rf_ram.memory\[562\]\[0\] _03860_ _03861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_41_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__14049__A1 mod.u_arbiter.i_wb_cpu_rdt\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14491__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07723__A1 _01857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_243_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_228_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08612_ mod.u_cpu.rf_ram.memory\[132\]\[1\] mod.u_cpu.rf_ram.memory\[133\]\[1\] mod.u_cpu.rf_ram.memory\[134\]\[1\]
+ mod.u_cpu.rf_ram.memory\[135\]\[1\] _01893_ _02054_ _02919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_209_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09592_ _03374_ _03720_ _03806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__13647__I1 mod.u_arbiter.i_wb_cpu_rdt\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08118__I3 mod.u_cpu.rf_ram.memory\[35\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08543_ _02216_ mod.u_cpu.rf_ram.memory\[294\]\[1\] _02849_ _01504_ _02850_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_82_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_224_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_208_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_243_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_211_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08474_ _01729_ _02780_ _02781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_196_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_210_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_211_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07425_ _01728_ mod.u_cpu.rf_ram.memory\[406\]\[0\] _01731_ _01732_ _01733_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_196_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09228__A1 _03485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_143_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11035__A1 _04821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12083__I0 _05533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_183_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07356_ _01663_ _01664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_17_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12783__A1 _05649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11830__I0 _05364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07287_ _01573_ _01594_ _01595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10633__I1 _04532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_40_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_191_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09026_ _03315_ _03327_ _03328_ _03330_ _01394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_156_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13732__B1 _06737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09400__A1 _03635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07637__S1 _01932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_176_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09951__A2 _03722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14834__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07962__A1 _02245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09928_ _04054_ mod.u_cpu.rf_ram.memory\[52\]\[1\] _04059_ _04061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_63_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08301__B _02102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09703__A2 _03892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_258_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09859_ _03809_ _04013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_74_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07565__I1 mod.u_cpu.rf_ram.memory\[369\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_234_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12870_ _06069_ _01104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__14984__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_233_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11649__I0 _05222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_227_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11821_ _05239_ _03829_ _05359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_3179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_215_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13263__A2 _06360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_214_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14540_ _00394_ net3 mod.u_cpu.rf_ram.memory\[417\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_202_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_11752_ _03884_ _05312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_14_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_215_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_214_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10321__I0 _04330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10703_ _04596_ _00410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_14471_ _00325_ net3 mod.u_cpu.rf_ram.memory\[452\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12049__I _03770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14212__A1 _03968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11683_ _05132_ _05265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08690__A2 _02993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_197_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11026__A1 _04412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13422_ _03377_ _03668_ net5 _06509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__12074__I0 _05521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10634_ _04550_ _00387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_10_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_259_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08690__C _02660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_167_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13353_ _06448_ _06449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_127_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10565_ _04369_ _04447_ _04503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__14364__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12304_ _05679_ mod.u_cpu.rf_ram.memory\[186\]\[0\] _05687_ _05688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_13284_ _06368_ _06382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_154_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10496_ _04457_ _04443_ _04458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_120_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15023_ _00877_ net3 mod.u_cpu.rf_ram.memory\[205\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_68_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13869__A4 _06283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12235_ _05593_ _05640_ _05641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_108_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10001__A2 _04109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12166_ _04379_ _05319_ _05594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_39_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11117_ _04879_ _04880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_122_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_256_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12097_ _04965_ _05543_ _05547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07606__I _01850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09093__I _03297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtiny_user_project_50 io_out[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_209_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_61 io_out[17] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_5060 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11888__I0 _05406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11048_ _04831_ _04822_ _04832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xtiny_user_project_72 io_out[28] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_5071 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5082 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07705__A1 _01711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtiny_user_project_83 la_data_out[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_92_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5093 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xtiny_user_project_94 la_data_out[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_188_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07800__S1 _02107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09821__I _03984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14807_ _00661_ net3 mod.u_cpu.rf_ram.memory\[284\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10967__I _03884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12999_ _06161_ _06164_ _06169_ _01133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_3691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_233_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_205_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_14738_ _00592_ net3 mod.u_cpu.rf_ram.memory\[318\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09042__B _03345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_221_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_205_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_178_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08130__A1 _02156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2990 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_221_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_221_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14669_ _00523_ net3 mod.u_cpu.rf_ram.memory\[353\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_60_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08681__A2 mod.u_cpu.rf_ram.memory\[208\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07210_ _01515_ _01518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08190_ _02457_ _02497_ _02498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__14707__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07141_ _01449_ mod.u_cpu.cpu.immdec.imm19_12_20\[5\] _01450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__12765__A1 _03950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14174__I _03928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10408__S _04397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_238_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14857__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13190__A1 _06116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07974_ mod.u_cpu.rf_ram.memory\[96\]\[0\] mod.u_cpu.rf_ram.memory\[97\]\[0\] mod.u_cpu.rf_ram.memory\[98\]\[0\]
+ mod.u_cpu.rf_ram.memory\[99\]\[0\] _02125_ _02127_ _02282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_228_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_214_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09713_ _03901_ _00115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09932__S _04063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11879__I0 _05383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09644_ _03846_ _00101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_67_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_215_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09731__I _03738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14237__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09575_ _03740_ mod.u_cpu.rf_ram.memory\[571\]\[0\] _03792_ _03793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_43_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_231_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11256__A1 _04973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08526_ _01872_ _02825_ _02832_ _01887_ _02833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__08347__I _02218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08121__A1 _02329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_211_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_211_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08457_ _01660_ _02764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__14387__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_212_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07408_ _01527_ _01716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_184_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_211_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15632__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08388_ _02692_ mod.u_cpu.rf_ram.memory\[420\]\[1\] _02694_ _02695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_137_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07339_ _01646_ _01647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_109_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_192_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10350_ _04348_ mod.u_cpu.rf_ram.memory\[466\]\[0\] _04357_ _04358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_191_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_191_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09009_ _01430_ _03313_ _03260_ _03314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_118_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10281_ _04043_ _04311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_191_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12020_ _05484_ mod.u_cpu.rf_ram.memory\[214\]\[1\] _05495_ _05497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_105_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11031__I1 _04819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_215_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_238_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15012__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_265_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13971_ mod.u_arbiter.i_wb_cpu_rdt\[5\] _06940_ _06941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_47_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_219_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07538__I1 _01840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_219_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_207_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_189_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12922_ _06103_ _01122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_262_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_207_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08685__C _01489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_234_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15641_ _01412_ net3 mod.u_cpu.rf_ram.memory\[269\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_132_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15162__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12853_ _06056_ _06057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08750__I3 mod.u_cpu.rf_ram.memory\[107\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_261_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13163__I _06204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11804_ _05132_ _05348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15572_ _01343_ net3 mod.u_arbiter.i_wb_cpu_dbus_dat\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12295__I0 _05677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12784_ _06010_ mod.u_cpu.rf_ram.memory\[131\]\[0\] _06012_ _06013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_2275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11798__A2 _05335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_30_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14523_ _00377_ net3 mod.u_cpu.rf_ram.memory\[426\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11735_ _05299_ _00739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_199_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08663__A2 _02969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11612__S _05215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_175_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12047__I0 _05501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14454_ _00308_ net3 mod.u_cpu.rf_ram.memory\[460\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_230_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11666_ _03665_ _04224_ _05252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_128_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13405_ mod.u_cpu.cpu.immdec.imm30_25\[0\] _06413_ _06357_ _06499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_10617_ _03940_ _04539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_14385_ _00239_ net3 mod.u_cpu.rf_ram.memory\[495\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11597_ _05205_ _00695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_183_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09088__I mod.u_cpu.cpu.state.o_cnt_r\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13336_ _06423_ _06430_ _06432_ _06433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_155_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10548_ _04486_ mod.u_cpu.rf_ram.memory\[434\]\[0\] _04491_ _04492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_115_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13267_ _06329_ _06365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_170_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10479_ _04430_ mod.u_cpu.rf_ram.memory\[446\]\[1\] _04444_ _04446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_142_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15006_ _00860_ net3 mod.u_cpu.rf_ram.memory\[210\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__13172__A1 _06047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_237_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12218_ _05628_ _00893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_155_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11022__I1 mod.u_cpu.rf_ram.memory\[358\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13198_ _06301_ _06304_ _06305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_9_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12149_ _02181_ _05580_ _05582_ _00870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_155_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_257_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07336__I _01494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15505__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_266_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07690_ _01752_ _01998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10533__I0 _04481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09551__I _03695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08351__A1 _02085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_252_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_225_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11238__A1 _04821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12286__I0 _05662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08167__I _01702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09360_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[21\] _03602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_244_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_240_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09151__I0 mod.u_arbiter.i_wb_cpu_rdt\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07537__S0 _01843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_178_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08311_ _02611_ _02614_ _02617_ _01742_ _02618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__12986__A1 _06063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09291_ _03541_ _03543_ _03544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_60_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09199__S _03469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_221_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08242_ _02156_ _02550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_127_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_193_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12738__A1 _05843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08173_ _02479_ _02480_ _02481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_158_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_203_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11321__I _03821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07124_ mod.u_cpu.cpu.state.genblk1.misalign_trap_sync_r _01433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_174_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15035__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_248_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12910__A1 _04913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08590__A1 _02688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_247_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07957_ _02170_ _02257_ _02264_ _02168_ _02265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_130_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15185__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_229_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_244_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07888_ _01851_ _02196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07145__A2 _01453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08342__A1 _02220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09627_ _03833_ _00097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_243_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_216_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09558_ _03700_ _03743_ _03778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_19_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_197_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08509_ _02665_ _02808_ _02815_ _02677_ _02816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_52_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_196_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_1243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09489_ _01460_ _03374_ _03715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_141_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11520_ _05147_ mod.u_cpu.rf_ram.memory\[280\]\[1\] _05153_ _05155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_200_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_197_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_196_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_180_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_221_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11451_ _05105_ _05106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12327__I _05667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08026__B _02333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10402_ _04365_ mod.u_cpu.rf_ram.memory\[458\]\[0\] _04393_ _04394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_14170_ _06047_ _07078_ _01395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_11382_ _05050_ mod.u_cpu.rf_ram.memory\[302\]\[1\] _05059_ _05061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__13867__B _06791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_194_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13121_ _03774_ _06249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_152_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10333_ _04345_ mod.u_cpu.rf_ram.memory\[46\]\[1\] _04342_ _04346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_125_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09358__B1 _03555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11004__I1 _04661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13052_ _03923_ _06204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_219_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10264_ _04288_ mod.u_cpu.rf_ram.memory\[47\]\[1\] _04295_ _04297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_133_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15528__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14402__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12003_ _05485_ _00821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_121_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_239_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10195_ _04248_ _04249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_65_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10763__I0 _04626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_266_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13094__S _06231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11468__A1 _03993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13954_ _03441_ _06917_ _06918_ _06926_ _06927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_98_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10515__I0 _04469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14552__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08333__A1 _02197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07767__S0 _01925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_234_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_12905_ _05657_ _06092_ _06093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_62_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13209__A2 _06300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13885_ _06735_ _06672_ _06875_ _06876_ _06877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_59_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_263_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12268__I0 _05662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_185_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2050 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12836_ _06046_ _06047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_15624_ _01395_ net3 mod.u_cpu.cpu.state.genblk1.misalign_trap_sync_r vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2061 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_50_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2072 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2083 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_226_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__12968__A1 _06142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15555_ _01326_ net3 mod.u_cpu.cpu.branch_op vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2094 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10818__I1 mod.u_cpu.rf_ram.memory\[390\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12438__S _05777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12767_ _06001_ _01069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_203_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_203_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14506_ _00360_ net3 mod.u_cpu.rf_ram.memory\[434\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11718_ _05288_ _00733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_187_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15486_ _01257_ net3 mod.u_arbiter.i_wb_cpu_dbus_adr\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_187_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12698_ _05934_ mod.u_cpu.rf_ram.memory\[140\]\[0\] _05956_ _05957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_30_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14437_ _00291_ net3 mod.u_cpu.rf_ram.memory\[46\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11649_ _05222_ mod.u_cpu.rf_ram.memory\[24\]\[0\] _05240_ _05241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_128_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11141__I _04879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15058__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13393__A1 _06442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_200_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_190_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14368_ _00222_ net3 mod.u_cpu.rf_ram.memory\[503\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12440__I0 _05761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13319_ _06415_ _06416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10980__I _03903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_192_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14299_ _00153_ net3 mod.u_cpu.rf_ram.memory\[538\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_115_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09546__I _03701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_254_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_171_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13696__A2 _06306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08860_ _01468_ _03051_ _03166_ _03167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_97_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07811_ _02115_ mod.u_cpu.rf_ram.memory\[174\]\[0\] _02118_ _01771_ _02119_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_229_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08791_ mod.u_cpu.rf_ram.memory\[78\]\[1\] mod.u_cpu.rf_ram.memory\[79\]\[1\] _01517_
+ _03098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_81_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_211_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07742_ mod.u_cpu.rf_ram.memory\[144\]\[0\] mod.u_cpu.rf_ram.memory\[145\]\[0\] mod.u_cpu.rf_ram.memory\[146\]\[0\]
+ mod.u_cpu.rf_ram.memory\[147\]\[0\] _02048_ _02049_ _02050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__09281__I _03517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_253_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10131__A1 _04201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07673_ _01750_ _01981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_225_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09412_ _03439_ mod.u_scanchain_local.module_data_in\[65\] _03647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_92_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_241_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_206_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12959__A1 mod.u_arbiter.i_wb_cpu_ibus_adr\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09343_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[18\] _03588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_80_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_209_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13620__A2 _04989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_178_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_33_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11631__A1 _02012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09274_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[7\] _03529_ _03530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__10434__A2 _04413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_240_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_193_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_194_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08225_ _02532_ _02533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_193_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13384__A1 _03663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08156_ _02462_ _02463_ _02464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_174_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10198__A1 _04251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14425__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_174_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08087_ mod.u_cpu.rf_ram.memory\[29\]\[0\] _02395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_106_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13687__A2 _06485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_249_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_216_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_251_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10745__I0 _04622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14575__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08563__A1 _01697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_88_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4903 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4914 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08989_ _03267_ _03278_ _03293_ _03294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XTAP_4925 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4936 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13706__I _06669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4947 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_169_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4958 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_180_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__12498__I0 _05813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4969 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08315__A1 _02225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_216_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10951_ _04764_ _00490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_249_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_232_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_186_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10130__I _04142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_232_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_204_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13670_ _06651_ _06657_ _06681_ _01292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_73_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10882_ _04695_ mod.u_cpu.rf_ram.memory\[380\]\[0\] _04717_ _04718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_182_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_227_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_12621_ _05904_ mod.u_cpu.rf_ram.memory\[151\]\[0\] _05905_ _05906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_231_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_244_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09815__A1 _03757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_145_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13611__A2 _03687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_15340_ _01115_ net3 mod.u_cpu.rf_ram.memory\[96\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_200_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_196_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15200__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12552_ _05859_ _00996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_184_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_11503_ _04959_ _05143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_185_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_157_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15271_ _00028_ net4 mod.u_arbiter.i_wb_cpu_rdt\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_200_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12483_ _05815_ _00971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_184_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14222_ _00078_ net3 mod.u_cpu.rf_ram.memory\[9\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_8_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11434_ mod.u_cpu.rf_ram.memory\[293\]\[1\] _05065_ _05093_ _05095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_171_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11896__I _05309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15350__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_256_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14153_ _07066_ _01390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_125_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11365_ _05031_ _05050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_153_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10984__I0 _04772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13104_ _06238_ _01169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_125_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14918__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14175__I0 _07081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_180_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08270__I _02139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10316_ _04334_ _00285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_112_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14084_ _07021_ mod.u_cpu.rf_ram.memory\[113\]\[0\] _07022_ _07023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_11296_ _04999_ mod.u_cpu.rf_ram.memory\[316\]\[1\] _05001_ _05003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_4_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10305__I _04302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13035_ _05396_ _06193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11689__A1 _05139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10247_ _04125_ _04285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_105_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10736__I0 _04598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08554__A1 _01938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07988__S0 _02294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10178_ _04215_ mod.u_cpu.rf_ram.memory\[492\]\[1\] _04235_ _04237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_67_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_152_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12489__I0 _05807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14986_ _00840_ net3 mod.u_cpu.rf_ram.memory\[62\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08306__A1 _02593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_235_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_47_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13937_ _05792_ _06912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_207_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08857__A2 _03146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13850__A2 _06443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_262_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_13868_ _06365_ _06861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_223_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_15607_ _01378_ net3 mod.u_cpu.rf_ram.memory\[11\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12819_ _03751_ _05721_ _06036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_188_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13799_ _06339_ _06790_ _06796_ _06799_ _06800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__08609__A2 _02915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_210_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15538_ _01309_ net3 mod.u_cpu.cpu.immdec.imm24_20\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12661__I0 _05918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_241_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_241_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_187_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14448__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_176_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_15469_ _01243_ net3 mod.u_cpu.cpu.ctrl.o_ibus_adr\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_204_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_200_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_191_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_200_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12169__A2 _05595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13366__A1 _06326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08010_ _02303_ _02317_ _02318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_159_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12413__I0 _05761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_190_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_143_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14598__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08793__A1 _02161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_239_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09961_ _04083_ _00181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_143_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08912_ _02546_ mod.u_cpu.rf_ram.memory\[524\]\[1\] _03218_ _03219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__12716__I1 mod.u_cpu.rf_ram.memory\[138\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10215__I _04136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09892_ _04036_ mod.u_cpu.rf_ram.memory\[535\]\[1\] _04034_ _04037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_258_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08843_ _02191_ _03148_ _03149_ _02093_ _03150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_135_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11247__S _04966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08774_ _02477_ mod.u_cpu.rf_ram.memory\[116\]\[1\] _03080_ _03081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_100_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07524__I _01444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07725_ _01992_ _02021_ _02032_ _02007_ _02033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_72_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_214_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09896__I1 mod.u_cpu.rf_ram.memory\[534\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13841__A2 _06834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07656_ mod.u_cpu.rf_ram.memory\[301\]\[0\] _01964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__15223__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_213_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10885__I _04719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07587_ _01759_ _01894_ _01895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_240_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09326_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[15\] _03574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10407__A2 _04380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_178_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11604__A1 _03723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_181_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15373__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_194_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09257_ _03495_ _03516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_139_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_239_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08208_ _02483_ mod.u_cpu.rf_ram.memory\[566\]\[0\] _02514_ _02515_ _02516_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_154_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09188_ mod.u_arbiter.i_wb_cpu_rdt\[20\] mod.u_arbiter.i_wb_cpu_dbus_dat\[17\] _03464_
+ _03466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_153_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_193_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_182_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08459__S1 _01958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08139_ _01471_ _02382_ _02446_ _02447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_257_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11150_ _04758_ _04887_ _04902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_190_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10101_ _04180_ _04164_ _04181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_68_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_150_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11081_ _04855_ _00529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_5401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08536__A1 _02730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10032_ _04115_ mod.u_cpu.rf_ram.memory\[512\]\[1\] _04129_ _04131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_114_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_5434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_248_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_194_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_5456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13436__I _06510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14840_ _00694_ net3 mod.u_cpu.rf_ram.memory\[267\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_264_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07434__I _01741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_217_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14771_ _00625_ net3 mod.u_cpu.rf_ram.memory\[302\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11983_ _05470_ mod.u_cpu.rf_ram.memory\[216\]\[0\] _05472_ _05473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_84_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_263_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_244_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13832__A2 _03670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_264_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_13722_ _06463_ _06662_ _06729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08395__S0 _02688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10934_ _04752_ _00485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10646__A2 _04534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11843__A1 _04845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_260_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_205_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_232_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_182_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_220_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13653_ _06447_ _06660_ _06663_ _06664_ _06665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_44_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10865_ _01865_ _04705_ _04706_ _00462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_12604_ _05894_ _01013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__13596__A1 mod.u_arbiter.i_wb_cpu_dbus_adr\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_176_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_73_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13584_ _06612_ _01275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_197_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__09264__A2 _03521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10796_ _03924_ _04658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_197_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_15323_ _01101_ net3 mod.u_cpu.rf_ram_if.rdata0\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07275__A1 _01577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12535_ _05848_ _00990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_223_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_185_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_200_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14740__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13348__B2 _06401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15254_ _00010_ net4 mod.u_arbiter.i_wb_cpu_rdt\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_9_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12466_ _05789_ _05803_ _00966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09016__A2 mod.u_cpu.cpu.ctrl.i_iscomp vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13899__A2 _06140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_201_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14205_ _07076_ _07099_ _01410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_11417_ _05069_ mod.u_cpu.rf_ram.memory\[296\]\[1\] _05082_ _05084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_32_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15185_ _01038_ net3 mod.u_cpu.rf_ram.memory\[143\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_197_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_12397_ _05581_ _05750_ _05751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_99_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14136_ _07055_ mod.u_cpu.rf_ram.memory\[115\]\[1\] _07053_ _07056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_11348_ _04989_ _05038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_153_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08870__S1 _02473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_140_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14890__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14067_ _07010_ _07011_ _01359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_113_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11279_ _04852_ _04990_ _04991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10709__I0 _04598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09575__I0 _03740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13018_ _06181_ _03919_ _06182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08868__C _02555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13520__A1 mod.u_arbiter.i_wb_cpu_dbus_adr\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_95_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11382__I0 _05050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13346__I _06424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15246__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14969_ _00823_ net3 mod.u_cpu.rf_ram.memory\[575\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_82_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07510_ _01657_ _01818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_263_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11834__A1 _05367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08490_ _02664_ _02787_ _02796_ _02797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_63_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12882__I0 _06073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07502__A2 mod.u_cpu.rf_ram.memory\[446\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14270__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15396__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07441_ _01498_ _01749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_223_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_250_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_149_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_222_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08175__I _02175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12634__I0 _05907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07372_ _01679_ _01680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_176_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09111_ _03410_ mod.timer_irq _03411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08108__C _02415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_198_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13339__A1 _06434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09042_ _01432_ _03333_ _03345_ _03346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_148_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09007__A2 _03309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07947__C _02207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_175_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_191_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_198_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12011__A1 _04294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_198_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_209_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_172_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07519__I _01700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08081__I3 mod.u_cpu.rf_ram.memory\[15\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08861__S1 _02451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09944_ _04072_ _00175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_132_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_252_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09734__I _03917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09566__I0 _03764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08778__C _01717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13511__B2 _06566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09875_ _04024_ _04025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_219_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4007 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10176__I1 mod.u_cpu.rf_ram.memory\[492\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4018 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4029 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08826_ _02406_ _03132_ _03133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10876__A2 _04713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_246_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_79_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09670__S _03867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08757_ _02220_ _03063_ _03064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11125__I0 _04880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14613__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_245_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08794__B _03100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_226_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_214_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_199_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07708_ _01967_ _02015_ _02016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_38_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1904 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08688_ _02179_ mod.u_cpu.rf_ram.memory\[204\]\[1\] _02995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_96_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_199_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09494__A2 _01454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_242_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1926 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_202_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07639_ _01934_ _01946_ _01947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1948 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1959 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_110_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_241_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14763__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08085__I _02126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10650_ _04560_ mod.u_cpu.rf_ram.memory\[418\]\[1\] _04558_ _04561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_198_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_224_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09309_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[13\] mod.u_cpu.cpu.ctrl.o_ibus_adr\[12\] _03559_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07257__A1 _01505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11053__A2 _04822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15313__CLKN net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10581_ _04497_ _04514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_167_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12320_ _05692_ mod.u_cpu.rf_ram.memory\[189\]\[1\] _05697_ _05699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_182_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07857__C _02164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15119__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12251_ _05652_ _00902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_181_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13050__I0 _06199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10056__S _04149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_207_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11202_ _04936_ mod.u_cpu.rf_ram.memory\[330\]\[1\] _04934_ _04937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08757__A1 _02220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13750__A1 _03510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12553__A2 _05757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12182_ _05309_ _05604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_123_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_190_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11133_ _04014_ _04887_ _04891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_150_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15269__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08509__A1 _02665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11064_ _04842_ _00525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_62_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_49_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_249_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_49_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_101 la_data_out[19] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_153_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xtiny_user_project_112 la_data_out[30] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_10015_ _04120_ _00198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_5264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xtiny_user_project_123 la_data_out[41] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_5275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_209_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_134 la_data_out[52] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_92_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xtiny_user_project_145 la_data_out[63] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_64_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xtiny_user_project_156 wbs_dat_o[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_4552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_218_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14823_ _00677_ net3 mod.u_cpu.rf_ram.memory\[276\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__14293__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtiny_user_project_167 wbs_dat_o[17] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_76_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xtiny_user_project_178 wbs_dat_o[28] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_218_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_217_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13805__A2 _06452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_233_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11816__A1 _05355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_205_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14754_ _00608_ net3 mod.u_cpu.rf_ram.memory\[310\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_151_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11966_ _05450_ mod.u_cpu.rf_ram.memory\[539\]\[1\] _05459_ _05461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_3884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3895 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13705_ _06317_ _06644_ _06713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10917_ _03827_ _04741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_45_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07496__A1 _01802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14685_ _00539_ net3 mod.u_cpu.rf_ram.memory\[345\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_232_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11897_ _05412_ _05413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09312__C _03561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_189_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_204_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_220_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13636_ _06412_ _06649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_34_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10848_ _04682_ mod.u_cpu.rf_ram.memory\[385\]\[1\] _04691_ _04693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_220_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_220_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13567_ mod.u_arbiter.i_wb_cpu_dbus_adr\[17\] mod.u_arbiter.i_wb_cpu_dbus_adr\[18\]
+ _06599_ _06603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_185_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10779_ _04647_ _00435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_121_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_201_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12518_ _05837_ mod.u_cpu.rf_ram.memory\[167\]\[1\] _05835_ _05838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_15306_ _00067_ net4 mod.u_scanchain_local.module_data_in\[63\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_157_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13498_ _06537_ _06557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_117_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_12449_ _05786_ _05787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_15237_ _01090_ net3 mod.u_cpu.rf_ram.memory\[125\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_154_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07339__I _01646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_176_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08748__A1 _02585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13785__B _06786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15168_ _01021_ net3 mod.u_cpu.rf_ram.memory\[150\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_141_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08879__B _02609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14119_ _07045_ _01377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_119_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07990_ _01744_ _02298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_15099_ _00953_ net3 mod.u_cpu.rf_ram.memory\[176\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_119_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_262_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11355__I0 _05028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14636__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_228_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09660_ _03855_ _03859_ _03860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_28_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_228_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14049__A2 _06998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07723__A2 mod.u_cpu.rf_ram.memory\[270\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08611_ _02074_ _02917_ _01662_ _02918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_83_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09591_ _03804_ _03805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_55_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_227_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11525__S _05156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08542_ _02091_ _02848_ _02849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_224_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14786__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07802__I _02109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_247_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07487__A1 _01728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08473_ mod.u_cpu.rf_ram.memory\[365\]\[1\] _02780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__11324__I _04541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_251_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07424_ _01614_ _01732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_223_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07239__A1 _01520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11035__A2 _04822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07355_ _01538_ _01663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12083__I1 mod.u_cpu.rf_ram.memory\[212\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_210_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_176_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13980__A1 mod.u_arbiter.i_wb_cpu_rdt\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12783__A2 _06011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_109_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_191_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07286_ mod.u_cpu.rf_ram.memory\[501\]\[0\] _01594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_163_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09025_ _01428_ _03328_ _03329_ _03330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_164_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08739__A1 _02043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15411__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11594__I0 _05199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_254_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08789__B _01534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10604__S _04529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_160_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09927_ _04060_ _00170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_172_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_98_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15561__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09858_ _04012_ _00149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_219_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08911__A1 _02509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08762__I1 mod.u_cpu.rf_ram.memory\[121\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08809_ _01483_ _03088_ _03115_ _03116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__13099__I0 _06230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_206_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09789_ _03960_ _03961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_3147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_234_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_227_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11820_ _05358_ _00765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13799__A1 _06339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07712__I _01993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11751_ _05310_ _05311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_54_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07478__A1 _01773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_214_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_183_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_202_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_187_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_202_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_187_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10702_ _04584_ mod.u_cpu.rf_ram.memory\[40\]\[0\] _04595_ _04596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_187_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14470_ _00324_ net3 mod.u_cpu.rf_ram.memory\[452\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_199_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11682_ _04700_ _05263_ _05264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_42_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14212__A2 _05120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_186_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_202_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13421_ _06508_ _01216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12223__A1 _05581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11026__A2 _04780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10633_ mod.u_cpu.rf_ram.memory\[421\]\[1\] _04532_ _04548_ _04550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_224_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09639__I _03842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14509__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08978__A1 _01430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13352_ _06316_ _06448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13971__A1 mod.u_arbiter.i_wb_cpu_rdt\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10564_ _04502_ _00365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_139_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_194_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12303_ _05452_ _05686_ _05687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_13283_ _06380_ _06381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_10495_ _03790_ _04457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_136_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15091__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15022_ _00876_ net3 mod.u_cpu.rf_ram.memory\[205\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_136_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12234_ _03727_ _04227_ _05640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_108_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13574__I1 mod.u_arbiter.i_wb_cpu_dbus_adr\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11585__I0 _05194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14659__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12165_ _03894_ _05593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_190_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11116_ _04795_ _04879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_151_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_235_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_12096_ _05546_ _00853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_49_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08211__C _02518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtiny_user_project_40 io_oeb[32] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_51 io_out[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_5050 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11047_ _03973_ _04831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_5061 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xtiny_user_project_62 io_out[18] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_73 io_out[29] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_92_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5072 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07705__A2 _02012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_84 la_data_out[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_65_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08902__A1 _02507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5083 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5094 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xtiny_user_project_95 la_data_out[13] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_237_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_209_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_264_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14806_ _00660_ net3 mod.u_cpu.rf_ram.memory\[284\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_4393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_149_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_206_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12998_ _06164_ _06168_ _06169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_3692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07469__A1 _01728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14737_ _00591_ net3 mod.u_cpu.rf_ram.memory\[31\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11949_ _05405_ _05450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_166_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_233_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2980 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08130__A2 mod.u_cpu.rf_ram.memory\[44\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2991 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_205_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14668_ _00522_ net3 mod.u_cpu.rf_ram.memory\[353\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_203_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12214__A1 _05355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13619_ _06635_ _01287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_14599_ _00453_ net3 mod.u_cpu.rf_ram.memory\[388\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_146_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08969__A1 _01421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09549__I _03770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_192_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15434__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07140_ _01448_ _01449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_125_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_125_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13714__A1 _03364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15584__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13190__A2 mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_236_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07973_ _02079_ _02147_ _01481_ _02280_ _02281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_87_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_228_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09712_ mod.u_cpu.rf_ram.memory\[557\]\[1\] _03735_ _03897_ _03901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_101_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09643_ _03832_ mod.u_cpu.rf_ram.memory\[564\]\[1\] _03844_ _03846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_83_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_256_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_228_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_209_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09574_ _03758_ _03791_ _03792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12828__I0 _06038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_208_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08525_ _01874_ _02828_ _02831_ _01884_ _02832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11256__A2 _04969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12453__A1 _03289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_196_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08121__A2 mod.u_cpu.rf_ram.memory\[36\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_196_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08752__S0 _02211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_212_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_196_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08456_ _02711_ _02761_ _02762_ _01698_ _02763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_23_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07407_ _01709_ mod.u_cpu.rf_ram.memory\[414\]\[0\] _01713_ _01714_ _01715_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_91_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08387_ _02532_ _02693_ _02694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13253__I0 _06351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_211_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07338_ _01645_ _01646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_136_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_192_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_192_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07632__A1 _01507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14801__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07269_ _01516_ _01577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_118_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_192_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_247_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09008_ mod.u_cpu.cpu.alu.cmp_r _03313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_191_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13556__I1 mod.u_arbiter.i_wb_cpu_dbus_adr\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10280_ _04307_ _04309_ _04310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_152_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10519__A1 _04251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11567__I0 _05178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_183_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_2_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12613__I _05373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_254_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09194__I _03451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14951__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_266_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11319__I0 _05014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11229__I _04107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09137__A1 mod.u_arbiter.i_wb_cpu_rdt\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13970_ _03412_ _03614_ _06940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_47_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07538__I2 _01842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09932__I0 _04051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_219_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12921_ _06088_ mod.u_cpu.rf_ram.memory\[379\]\[0\] _06102_ _06103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12692__A1 _04643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15307__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_207_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_246_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15640_ _01411_ net3 mod.u_cpu.cpu.state.stage_two_req vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12852_ _03398_ _06056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_132_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07442__I _01749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_262_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11803_ _04539_ _05279_ _05347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_27_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_221_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15571_ _01342_ net3 mod.u_arbiter.i_wb_cpu_dbus_dat\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12783_ _05649_ _06011_ _06012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_215_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_265_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_215_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_202_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11734_ _05287_ mod.u_cpu.rf_ram.memory\[241\]\[1\] _05297_ _05299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XPHY_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__15457__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14522_ _00376_ net3 mod.u_cpu.rf_ram.memory\[426\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14331__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_186_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_230_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_203_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_30_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_202_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11665_ _05251_ _00717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_202_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14453_ _00307_ net3 mod.u_cpu.rf_ram.memory\[461\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__13244__I0 _06276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_202_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10058__I0 _04140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13404_ _06483_ _06492_ _06497_ _06498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_10616_ _04538_ _00381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_155_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14384_ _00238_ net3 mod.u_cpu.rf_ram.memory\[495\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_70_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11596_ _05194_ mod.u_cpu.rf_ram.memory\[267\]\[1\] _05203_ _05205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_127_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_196_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14481__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13335_ _06431_ _06432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_41_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10547_ _04201_ _04487_ _04491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_183_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13266_ _06361_ _06364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_155_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10478_ _04445_ _00336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_124_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12217_ _05609_ mod.u_cpu.rf_ram.memory\[198\]\[1\] _05626_ _05628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_15005_ _00859_ net3 mod.u_cpu.rf_ram.memory\[68\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_124_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13197_ _06302_ _06303_ _06304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_233_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10230__I0 _04249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12148_ _05581_ _05580_ _05582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_110_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10930__A1 _04749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_256_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10043__I _04090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12079_ _03841_ _05535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_133_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08876__C _02487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09923__I0 _04054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_238_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_213_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_206_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_80_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13290__S _06122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_178_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08310_ _02198_ mod.u_cpu.rf_ram.memory\[478\]\[1\] _02616_ _01751_ _02617_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__07537__S1 _01844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09290_ _03542_ _03538_ _03543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__12986__A2 _03335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_221_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_221_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08241_ _02546_ mod.u_cpu.rf_ram.memory\[524\]\[0\] _02548_ _02549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__14824__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10049__I0 _04117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_193_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08172_ mod.u_cpu.rf_ram.memory\[557\]\[0\] _02480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_165_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08183__I _02321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09064__B1 _03355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09603__A2 _03805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_158_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07123_ mod.u_cpu.cpu.decode.co_ebreak _01427_ _01424_ _01431_ _01432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XANTENNA__07614__A1 _01920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__14974__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11549__I0 _05162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07955__C _02252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12210__I1 _05622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_217_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_88_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10221__I0 _04267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_82_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12910__A2 _04570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_101_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07956_ _02174_ _02260_ _02263_ _01766_ _02264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_229_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_249_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_262_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07887_ _02188_ _02189_ _02194_ _01833_ _02195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__12674__A1 _04913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_210_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_46_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_228_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08342__A2 _02648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09626_ _03832_ mod.u_cpu.rf_ram.memory\[566\]\[1\] _03830_ _03833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__14354__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07262__I _01569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_216_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_244_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09557_ _03777_ _00083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_71_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_231_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_203_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12809__S _06027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08508_ _02668_ _02811_ _02814_ _01687_ _02815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_180_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09488_ _03713_ _03714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_51_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_197_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08439_ _01770_ _02745_ _02746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_145_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10329__S _04342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_200_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_200_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_197_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_260_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11450_ _03732_ _05105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_165_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08026__C _02291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10401_ _04242_ _04373_ _04393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11381_ _05060_ _00624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_164_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13867__C _06131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_180_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13120_ _03941_ _04708_ _06248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_125_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10332_ _04344_ _04345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_139_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09358__A1 _03554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13051_ _06203_ _01151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08405__I0 mod.u_cpu.rf_ram.memory\[440\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10263_ _02439_ _04295_ _04296_ _00270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_87_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12201__I1 _05617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_3_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12002_ _05484_ mod.u_cpu.rf_ram.memory\[215\]\[1\] _05481_ _05485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07437__I _01744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10212__I0 _04245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10194_ _04247_ _04248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07464__S0 _01753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_238_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10912__A1 _04611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10763__I1 mod.u_cpu.rf_ram.memory\[3\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09905__I0 _04036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13953_ _06920_ _05793_ _06925_ _06926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__08333__A2 _02639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_189_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07767__S1 _02071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12904_ _05720_ _06092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_228_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13884_ _06492_ _06311_ _06876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_98_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_261_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_250_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2040 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15623_ _01394_ net3 mod.u_cpu.cpu.mem_if.signbit vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__14847__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_185_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2051 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12835_ net5 _06046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_15_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2062 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2073 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2084 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15554_ _01325_ net3 mod.u_arbiter.i_wb_cpu_dbus_we vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2095 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12766_ _05992_ mod.u_cpu.rf_ram.memory\[134\]\[0\] _06000_ _06001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_163_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_99_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14505_ _00359_ net3 mod.u_cpu.rf_ram.memory\[435\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11717_ _05287_ mod.u_cpu.rf_ram.memory\[248\]\[1\] _05285_ _05288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10239__S _04278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12697_ _03904_ _05940_ _05956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_15485_ _01256_ net3 mod.u_arbiter.i_wb_cpu_dbus_adr\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11422__I _05031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_175_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14997__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11648_ _05239_ _03805_ _05240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_14436_ _00290_ net3 mod.u_cpu.rf_ram.memory\[46\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_204_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09597__A1 _03805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_174_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13393__A2 _06398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10038__I _04135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11579_ _05177_ _05194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_14367_ _00221_ net3 mod.u_cpu.rf_ram.memory\[504\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12440__I1 mod.u_cpu.rf_ram.memory\[172\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10451__I0 _04410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13318_ _06138_ _06415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_115_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14227__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_192_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_155_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14298_ _00152_ net3 mod.u_cpu.rf_ram.memory\[538\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_182_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_192_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13249_ _06276_ mod.u_cpu.rf_ram.memory\[92\]\[1\] _06348_ _06350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_124_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_35_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_257_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07810_ _02116_ _02117_ _02118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_97_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14377__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08790_ _03090_ _03092_ _03094_ _03096_ _03097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__10702__S _04595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09562__I _03781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15622__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07741_ _02042_ _02049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_244_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11703__I0 _05271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13853__B1 _06837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_226_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07672_ mod.u_cpu.rf_ram.memory\[272\]\[0\] mod.u_cpu.rf_ram.memory\[273\]\[0\] mod.u_cpu.rf_ram.memory\[274\]\[0\]
+ mod.u_cpu.rf_ram.memory\[275\]\[0\] _01957_ _01958_ _01980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_53_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10131__A2 _04202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_129_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09411_ mod.u_arbiter.i_wb_cpu_dbus_adr\[28\] _03561_ _03644_ _03645_ _03646_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_226_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12408__A1 _05187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_240_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_179_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09342_ _03568_ _03584_ _03586_ _03587_ _00058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_80_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08088__A1 _02369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12959__A2 _05783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_221_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09273_ _03524_ _03525_ _03529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_205_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_166_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15002__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13908__A1 _03681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08224_ _01635_ _02532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_138_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08155_ mod.u_cpu.rf_ram.memory\[551\]\[0\] _02463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_14_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_162_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10198__A2 _03873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08086_ mod.u_cpu.rf_ram.memory\[24\]\[0\] mod.u_cpu.rf_ram.memory\[25\]\[0\] mod.u_cpu.rf_ram.memory\[26\]\[0\]
+ mod.u_cpu.rf_ram.memory\[27\]\[0\] _02349_ _02393_ _02394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__08260__A1 _02566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15152__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12195__I0 _05609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08012__A1 _02283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_130_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08797__B _01618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_5627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08563__A2 mod.u_cpu.rf_ram.memory\[310\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09760__A1 _03747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_102_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4904 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4915 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09472__I _03697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08988_ _03279_ _03292_ _03256_ _03293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_4926 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_102_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4937 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_180_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4948 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07939_ _02245_ _02246_ _02247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_263_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4959 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_169_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10950_ _04753_ mod.u_cpu.rf_ram.memory\[36\]\[0\] _04763_ _04764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_243_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_232_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09609_ _03707_ _03748_ _03819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_44_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10881_ _04315_ _04709_ _04717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12539__S _05849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_12620_ _03879_ _05900_ _05905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_43_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_227_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__09815__A2 _03980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_71_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_12551_ _05858_ mod.u_cpu.rf_ram.memory\[163\]\[1\] _05856_ _05859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XPHY_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_145_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_237_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_106_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_185_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08037__B _01534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_11502_ _05142_ _00663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_200_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_157_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15270_ _00027_ net4 mod.u_arbiter.i_wb_cpu_rdt\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12482_ _05813_ mod.u_cpu.rf_ram.memory\[449\]\[0\] _05814_ _05815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_184_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_14221_ _07108_ _01417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_172_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11433_ _01946_ _05093_ _05094_ _00642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_184_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11386__A1 _04817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14152_ _07055_ mod.u_cpu.rf_ram.memory\[247\]\[1\] _07064_ _07066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_11364_ _05049_ _00618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_152_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13103_ _06237_ mod.u_cpu.rf_ram.memory\[102\]\[1\] _06234_ _06238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_10315_ _04330_ mod.u_cpu.rf_ram.memory\[472\]\[1\] _04332_ _04334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_98_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14083_ _03865_ _07014_ _07022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_98_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14175__I1 mod.u_cpu.rf_ram.memory\[88\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_193_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11295_ _05002_ _00596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11138__A1 _04749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_234_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12186__I0 _05605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15645__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_180_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13034_ _06192_ _01145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08003__A1 _02105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10246_ _04284_ _00265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_156_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_239_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08554__A2 mod.u_cpu.rf_ram.memory\[318\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09751__A1 _03711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07988__S1 _02295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_266_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10177_ _04236_ _00244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_67_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10522__S _04473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_255_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_226_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_266_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14985_ _00839_ net3 mod.u_cpu.rf_ram.memory\[61\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_93_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09503__A1 _03714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_235_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13936_ _06910_ _06911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11310__A1 _04873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_170_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_235_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_208_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13850__A3 _06466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_223_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13867_ _06823_ _06449_ _06791_ _06131_ _06860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_35_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_222_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15025__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15606_ _01377_ net3 mod.u_cpu.rf_ram.memory\[11\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12818_ _05962_ _06035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07630__I _01825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13798_ _06401_ _06798_ _06409_ _06799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_31_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12248__I _05432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15537_ _01308_ net3 mod.u_cpu.cpu.immdec.imm24_20\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12749_ _05843_ _05989_ _05990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_163_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__14012__B1 _06971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08490__A1 _02664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07293__A2 _01593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15468_ _01242_ net3 mod.u_cpu.cpu.ctrl.o_ibus_adr\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__15175__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_198_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13366__A2 _06391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14419_ _00273_ net3 mod.u_cpu.rf_ram.memory\[478\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_200_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_191_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15399_ _01174_ net3 mod.u_cpu.rf_ram.memory\[0\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_129_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_200_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_144_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08793__A2 mod.u_cpu.rf_ram.memory\[76\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_170_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09960_ _04071_ mod.u_cpu.rf_ram.memory\[524\]\[1\] _04081_ _04083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_170_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08911_ _02509_ _03217_ _03218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09891_ _04017_ _04036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08842_ _02272_ mod.u_cpu.rf_ram.memory\[44\]\[1\] _03149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_111_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08773_ _01682_ _03079_ _03080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_245_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_211_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07724_ _01997_ _02025_ _02031_ _02005_ _02032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__08928__S0 _02528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_225_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_214_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07655_ _01644_ _01963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_26_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_53_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_241_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_198_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13542__I _06583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_198_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07586_ mod.u_cpu.rf_ram.memory\[365\]\[0\] _01894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_25_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13054__A1 _03858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07540__I _01457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09325_ _03568_ _03572_ _03573_ _00055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__15518__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12158__I _03712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11604__A2 _04779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12801__A1 _03985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_222_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_167_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_194_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_139_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09256_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[4\] _03514_ _03515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_103_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08207_ _02306_ _02515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_21_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13357__A2 _06451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09187_ _03465_ _00022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_166_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13601__I0 mod.u_cpu.rf_ram.memory\[329\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11368__A1 _04766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__14542__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08138_ _01475_ _02419_ _02445_ _02446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__08233__A1 _02523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_179_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09430__B1 _03493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10040__A1 _03991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09981__A1 _03933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_253_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08069_ _01551_ _02377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10406__I _03924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_255_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10100_ _03828_ _04180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_161_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11080_ _04841_ mod.u_cpu.rf_ram.memory\[350\]\[1\] _04853_ _04855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_108_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_249_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_216_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__12868__A1 _05896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14692__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08536__A2 _02842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09733__A1 _03711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10031_ _04130_ _00204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_5424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_237_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11540__A1 _04749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_130_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_208_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_217_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08919__S0 _02560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15048__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10141__I _03872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14770_ _00624_ net3 mod.u_cpu.rf_ram.memory\[302\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_4789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11982_ _05283_ _05471_ _05472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_90_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09930__I _04002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_186_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13721_ _06717_ _06727_ _06475_ _06728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__08395__S1 _02475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10933_ _04739_ mod.u_cpu.rf_ram.memory\[372\]\[1\] _04750_ _04752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_90_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_204_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11843__A2 _05374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_205_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13652_ _06129_ _06664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_10864_ _04611_ _04705_ _04706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_231_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__14093__I0 _07028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_220_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07450__I _01757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15198__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12603_ _05887_ mod.u_cpu.rf_ram.memory\[154\]\[0\] _05893_ _05894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_73_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_213_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13596__A2 _03694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_197_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10795_ _04657_ _00441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_13583_ mod.u_arbiter.i_wb_cpu_dbus_adr\[24\] mod.u_arbiter.i_wb_cpu_dbus_adr\[25\]
+ _06609_ _06612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XPHY_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__11901__S _05414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_262_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_200_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15322_ _01100_ net3 mod.u_cpu.rf_ram_if.rgnt vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_160_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07275__A2 mod.u_cpu.rf_ram.memory\[470\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12534_ mod.u_cpu.rf_ram.memory\[429\]\[1\] _05765_ _05846_ _05848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_157_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_184_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_200_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13401__B _06494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15253_ _00009_ net4 mod.u_arbiter.i_wb_cpu_rdt\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_8_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12465_ _01433_ _03284_ _03377_ _05802_ _05803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_201_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14204_ _06153_ _07098_ _07099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_11416_ _05083_ _00636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_165_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12396_ _04700_ _04335_ _05750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_15184_ _01037_ net3 mod.u_cpu.rf_ram.memory\[143\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_153_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11347_ _03849_ _05037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_14135_ _06903_ _07055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_119_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_119_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11278_ _04989_ _04990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_14066_ mod.u_arbiter.i_wb_cpu_rdt\[30\] _06937_ _07004_ mod.u_arbiter.i_wb_cpu_dbus_dat\[30\]
+ _07011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__12859__A1 mod.u_cpu.rf_ram_if.rtrig1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10709__I1 mod.u_cpu.rf_ram.memory\[408\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__13627__I _06415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13017_ _04982_ _06181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_10229_ _04272_ _04263_ _04273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13520__A2 _03669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10252__S _04286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_230_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_227_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__13808__B1 _06807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_208_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_254_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_208_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14968_ _00822_ net3 mod.u_cpu.rf_ram.memory\[575\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_66_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__12331__I0 _05692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_207_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_223_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_223_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13919_ _03403_ _06649_ _06896_ _06897_ _06898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__14415__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11834__A2 _05335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14899_ _00753_ net3 mod.u_cpu.rf_ram.memory\[235\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__13362__I _06391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11083__S _04856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_223_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07440_ mod.u_cpu.rf_ram.memory\[416\]\[0\] mod.u_cpu.rf_ram.memory\[417\]\[0\] mod.u_cpu.rf_ram.memory\[418\]\[0\]
+ mod.u_cpu.rf_ram.memory\[419\]\[0\] _01745_ _01747_ _01748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_90_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13036__A1 _05732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14084__I0 _07021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_223_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07371_ _01660_ _01679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_206_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_149_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12634__I1 mod.u_cpu.rf_ram.memory\[14\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_241_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11598__A1 _04792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11811__S _05352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09255__A3 _03503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09110_ _03409_ _03410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__14565__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_175_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08463__A1 _01858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09041_ _03336_ _03341_ _03344_ mod.u_cpu.cpu.genblk3.csr.mstatus_mie _03345_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_129_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11610__I _05119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_198_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_191_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12011__A2 _04026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08124__C _01828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_239_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09943_ _04071_ mod.u_cpu.rf_ram.memory\[527\]\[1\] _04069_ _04072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_217_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_131_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_258_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09715__A1 _03870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_225_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09874_ _03768_ _03786_ _04024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11522__A1 _05110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4008 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07535__I _01825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4019 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08825_ mod.u_cpu.rf_ram.memory\[21\]\[1\] _03132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_100_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08756_ mod.u_cpu.rf_ram.memory\[103\]\[1\] _03063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_72_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08794__C _02086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07707_ mod.u_cpu.rf_ram.memory\[263\]\[0\] _02015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_2_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08687_ mod.u_cpu.rf_ram.memory\[205\]\[1\] _02994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_54_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1905 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15340__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1927 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14908__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07638_ mod.u_cpu.rf_ram.memory\[293\]\[0\] _01946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1938 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_214_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_213_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07270__I _01560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1949 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14075__I0 _06904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_214_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_202_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_110_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07569_ _01759_ _01876_ _01877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_179_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11721__S _05290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_224_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09308_ _03552_ _03547_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[10\] _03543_ _03558_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__10636__I0 _04523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15490__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10580_ _04513_ _00370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_110_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10261__A1 _04294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09239_ _03499_ _03500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_155_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12389__I0 _05745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12250_ _05645_ mod.u_cpu.rf_ram.memory\[195\]\[0\] _05651_ _05652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_182_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_257_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_266_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11201_ _04879_ _04936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_163_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10013__A1 _03969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12181_ _05603_ _00881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13750__A2 mod.u_arbiter.i_wb_cpu_rdt\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11132_ _04890_ _00545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_123_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13447__I _06513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08509__A2 _02808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11063_ _04841_ mod.u_cpu.rf_ram.memory\[352\]\[1\] _04839_ _04842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07445__I _01752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xtiny_user_project_102 la_data_out[20] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_77_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10014_ _04117_ mod.u_cpu.rf_ram.memory\[515\]\[0\] _04119_ _04120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_5254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_231_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13891__B _06800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtiny_user_project_113 la_data_out[31] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_5265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xtiny_user_project_124 la_data_out[42] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_231_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14438__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_209_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_188_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_264_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xtiny_user_project_135 la_data_out[53] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_5287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_237_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xtiny_user_project_146 user_irq[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_4542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14822_ _00676_ net3 mod.u_cpu.rf_ram.memory\[276\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_4553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xtiny_user_project_157 wbs_dat_o[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_236_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xtiny_user_project_168 wbs_dat_o[18] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_179 wbs_dat_o[29] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_4575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_149_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_4597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_264_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_14753_ _00607_ net3 mod.u_cpu.rf_ram.memory\[311\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11816__A2 _05335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11965_ _05460_ _00808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3896 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_260_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_205_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13704_ _06470_ _06711_ _06480_ _06320_ _06712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_60_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14588__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10916_ _04740_ _00479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_229_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14684_ _00538_ net3 mod.u_cpu.rf_ram.memory\[345\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_60_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11896_ _05309_ _05412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07180__I _01487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08209__C _02489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13635_ _06642_ _06645_ _06646_ _06647_ _06648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_73_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10847_ _04692_ _00458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_125_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_201_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_13566_ _06602_ _01267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_160_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10778_ mod.u_cpu.rf_ram.memory\[397\]\[1\] _04532_ _04645_ _04647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_160_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08835__I3 mod.u_cpu.rf_ram.memory\[55\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15305_ _00066_ net4 mod.u_scanchain_local.module_data_in\[62\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_185_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08996__A2 mod.u_cpu.cpu.bufreg.i_sh_signed vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12517_ _05806_ _05837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_118_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_199_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13497_ _06556_ _01244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_117_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15236_ _01089_ net3 mod.u_cpu.rf_ram.memory\[125\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_161_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12448_ mod.u_arbiter.i_wb_cpu_ibus_adr\[1\] _05784_ _05785_ _05786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_126_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10046__I _04135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15167_ _01020_ net3 mod.u_cpu.rf_ram.memory\[151\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12379_ _05293_ _05726_ _05739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_181_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15213__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_236_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14118_ _07043_ mod.u_cpu.rf_ram.memory\[11\]\[0\] _07044_ _07045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_158_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15098_ _00952_ net3 mod.u_cpu.rf_ram.memory\[176\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_113_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14049_ mod.u_arbiter.i_wb_cpu_rdt\[25\] _06998_ _06993_ mod.u_arbiter.i_wb_cpu_dbus_dat\[25\]
+ _06999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_80_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_140_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07355__I _01538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input2_I io_in[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__15363__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08610_ mod.u_cpu.rf_ram.memory\[144\]\[1\] mod.u_cpu.rf_ram.memory\[145\]\[1\] mod.u_cpu.rf_ram.memory\[146\]\[1\]
+ mod.u_cpu.rf_ram.memory\[147\]\[1\] _02085_ _02049_ _02917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_09590_ _03803_ _03804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_255_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12304__I0 _05679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_209_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08541_ mod.u_cpu.rf_ram.memory\[295\]\[1\] _02848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_165_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13092__I _06204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_247_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08472_ mod.u_cpu.rf_ram.memory\[360\]\[1\] mod.u_cpu.rf_ram.memory\[361\]\[1\] mod.u_cpu.rf_ram.memory\[362\]\[1\]
+ mod.u_cpu.rf_ram.memory\[363\]\[1\] _02751_ _02748_ _02779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__08186__I _01705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10866__I0 _04698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08684__A1 _02230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07487__A2 mod.u_cpu.rf_ram.memory\[436\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_250_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_165_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07423_ _01729_ _01730_ _01731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_168_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_206_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07354_ _01661_ _01662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_148_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_13_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11291__I0 _04999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13980__A2 _06938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07285_ mod.u_cpu.rf_ram.memory\[496\]\[0\] mod.u_cpu.rf_ram.memory\[497\]\[0\] mod.u_cpu.rf_ram.memory\[498\]\[0\]
+ mod.u_cpu.rf_ram.memory\[499\]\[0\] _01540_ _01570_ _01593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_164_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_191_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09024_ mod.u_arbiter.i_wb_cpu_dbus_dat\[0\] mod.u_arbiter.i_wb_cpu_dbus_dat\[16\]
+ mod.u_arbiter.i_wb_cpu_dbus_dat\[8\] mod.u_arbiter.i_wb_cpu_dbus_dat\[24\] mod.u_cpu.cpu.bufreg.lsb\[1\]
+ mod.u_cpu.cpu.bufreg.lsb\[0\] _03329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_164_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09936__A1 _03818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13732__A2 _06657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12372__S _05733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_254_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_144_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__13267__I _06329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_259_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09926_ _04051_ mod.u_cpu.rf_ram.memory\[52\]\[0\] _04059_ _04060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_132_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13496__A1 _03635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09681__S _03874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07265__I _01510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09857_ _03999_ mod.u_cpu.rf_ram.memory\[540\]\[1\] _04010_ _04012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_246_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_213_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_218_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08808_ _02337_ _03097_ _03114_ _02380_ _03115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_3115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08762__I2 mod.u_cpu.rf_ram.memory\[122\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14730__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09788_ _03959_ _03960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08739_ _02043_ _03042_ _03045_ _01695_ _03046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__13799__A2 _06790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_227_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_199_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_242_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_199_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11750_ _05309_ _05310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_199_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_199_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10482__A1 _04307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_35 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10701_ _04511_ _03933_ _04595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_241_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14880__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11681_ _05262_ _05263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_230_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_198_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13420_ _06354_ mod.u_cpu.rf_ram.memory\[339\]\[1\] _06506_ _06508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_186_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10632_ _01754_ _04548_ _04549_ _00386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__12223__A2 _05632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11282__I0 _04976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_220_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13351_ _06441_ _06390_ _06447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_139_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10563_ _04498_ mod.u_cpu.rf_ram.memory\[432\]\[1\] _04500_ _04502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08978__A2 mod.u_arbiter.i_wb_cpu_dbus_dat\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_210_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13971__A2 _06940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11982__A1 _05283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15236__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12302_ _05667_ _05686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_155_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14220__I0 _03735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13282_ _06328_ _06379_ _06380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_143_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10494_ _04456_ _00341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_15021_ _00875_ net3 mod.u_cpu.rf_ram.memory\[73\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12233_ _05639_ _00897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13723__A2 _06668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_194_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09655__I _03757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12164_ _05592_ _00875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_155_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14260__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15386__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11115_ _04878_ _00540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_155_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12095_ _05533_ mod.u_cpu.rf_ram.memory\[66\]\[1\] _05544_ _05546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_96_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07175__I _01482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_249_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xtiny_user_project_30 io_oeb[22] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_11046_ _04830_ _00519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xtiny_user_project_41 io_oeb[33] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_5040 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xtiny_user_project_52 io_out[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_5051 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xtiny_user_project_63 io_out[19] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_5062 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xtiny_user_project_74 io_out[30] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_265_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5073 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5084 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xtiny_user_project_85 la_data_out[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_4350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_96 la_data_out[14] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_37_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5095 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_237_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_225_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_4361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14805_ _00659_ net3 mod.u_cpu.rf_ram.memory\[285\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_4394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11425__I _04995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12997_ _06166_ _03404_ _06167_ _05780_ _03373_ _06168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_188_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10848__I0 _04682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14736_ _00590_ net3 mod.u_cpu.rf_ram.memory\[31\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11948_ _02407_ _05447_ _05449_ _00802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__07469__A2 mod.u_cpu.rf_ram.memory\[428\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2970 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12462__A2 _03406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_232_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2981 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_205_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_205_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2992 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14667_ _00521_ net3 mod.u_cpu.rf_ram.memory\[354\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_127_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11879_ _05383_ mod.u_cpu.rf_ram.memory\[71\]\[1\] _05398_ _05400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_127_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_242_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_220_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13618_ _06581_ mod.u_cpu.rf_ram.memory\[319\]\[1\] _06633_ _06635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08418__A1 _02526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12214__A2 _05611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14598_ _00452_ net3 mod.u_cpu.rf_ram.memory\[388\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08969__A2 mod.u_cpu.cpu.branch_op vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13549_ mod.u_arbiter.i_wb_cpu_dbus_adr\[9\] mod.u_arbiter.i_wb_cpu_dbus_adr\[10\]
+ _06589_ _06593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_185_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_145_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_161_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14603__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_195_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15219_ _01072_ net3 mod.u_cpu.rf_ram.memory\[133\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__13714__A2 _06657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08402__C _01979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07972_ _02148_ _02232_ _02279_ _02280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__14753__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09711_ _02480_ _03897_ _03900_ _00114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_68_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_214_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_228_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07157__A1 _01464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13815__I _06431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09642_ _03845_ _00100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_68_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15109__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09573_ _03790_ _03791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_83_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08524_ _01879_ mod.u_cpu.rf_ram.memory\[342\]\[1\] _02830_ _01867_ _02831_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_36_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13650__A1 _06320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_212_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_251_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_169_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_224_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08752__S1 _02386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08455_ _01496_ mod.u_cpu.rf_ram.memory\[380\]\[1\] _02762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_223_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_212_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__15259__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07406_ _01524_ _01714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_17_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08386_ mod.u_cpu.rf_ram.memory\[421\]\[1\] _02693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_211_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13402__A1 _06381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_260_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10216__A1 _04262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11264__I0 _04978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07337_ _01644_ _01645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_177_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11070__I _04847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_129_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07268_ _01556_ mod.u_cpu.rf_ram.memory\[468\]\[0\] _01575_ _01576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__14283__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11016__I0 _04803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09007_ _03308_ _03309_ _03312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_3_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13705__A2 _06644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07199_ _01506_ _01507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_118_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_145_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10519__A2 _03911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08312__C _01678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_263_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_266_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09137__A2 _03410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09909_ _04048_ _00164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_150_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12141__A1 _04930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_247_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12920_ _05888_ _04704_ _06102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_115_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07538__I3 _01845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12692__A2 _05952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12851_ _06052_ _06055_ _01099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_2211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11802_ _05346_ _00759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15570_ _01341_ net3 mod.u_arbiter.i_wb_cpu_dbus_dat\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09696__I0 _03877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13641__A1 _03297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12782_ _05919_ _06011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_214_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_14521_ _00375_ net3 mod.u_cpu.rf_ram.memory\[427\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11733_ _05298_ _00738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_199_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_203_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_261_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_199_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_203_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14452_ _00306_ net3 mod.u_cpu.rf_ram.memory\[461\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_109_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11664_ _05250_ mod.u_cpu.rf_ram.memory\[257\]\[1\] _05247_ _05251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_230_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13403_ _06432_ _06403_ _06496_ _06497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__14626__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_168_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10615_ _04537_ mod.u_cpu.rf_ram.memory\[424\]\[1\] _04535_ _04538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_128_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14383_ _00237_ net3 mod.u_cpu.rf_ram.memory\[496\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09073__A1 _03371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11595_ _05204_ _00694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_155_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13334_ _06133_ _06431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_128_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07623__A2 _01917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08820__A1 _02411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10546_ _04490_ _00359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_109_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_259_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13265_ _06362_ _06363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_157_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10477_ _04423_ mod.u_cpu.rf_ram.memory\[446\]\[0\] _04444_ _04445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_6_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09385__I _03563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15004_ _00858_ net3 mod.u_cpu.rf_ram.memory\[68\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__14776__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12755__I0 _05992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12216_ _05627_ _00892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_170_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_237_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13196_ _05782_ mod.u_arbiter.i_wb_cpu_rdt\[13\] _06303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_97_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10230__I1 mod.u_cpu.rf_ram.memory\[484\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12147_ _05487_ _05581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_151_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12078_ _05534_ _00847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_81_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11029_ _01903_ _04816_ _04818_ _00514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_65_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08887__A1 _02455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_264_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_266_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09687__I0 _03877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15401__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_252_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_233_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_233_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14719_ _00573_ net3 mod.u_cpu.rf_ram.memory\[328\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_244_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_205_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07311__A1 _01602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08240_ _02509_ _02547_ _02548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_75_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_221_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_203_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08171_ _01925_ _02479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_14_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__10049__I1 mod.u_cpu.rf_ram.memory\[510\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_192_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15551__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09064__A1 _03362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09064__B2 _03364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07122_ _01428_ _01429_ _01430_ _01431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_174_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10435__S _04413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13699__A1 _03364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12746__I0 _05984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09295__I mod.u_cpu.cpu.ctrl.o_ibus_adr\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07808__I _01862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_173_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10221__I1 mod.u_cpu.rf_ram.memory\[486\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10234__I _04248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09119__A2 _03392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07955_ _02249_ mod.u_cpu.rf_ram.memory\[246\]\[0\] _02262_ _02252_ _02263_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_102_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_229_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_214_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_233_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08878__A1 _02592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08639__I mod.u_cpu.rf_ram.memory\[173\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07886_ _02191_ _02192_ _02193_ _01666_ _02194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__13871__A1 _06840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_256_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07543__I _01850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09625_ _03763_ _03832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10685__A1 _04315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_216_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_216_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11065__I _04802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13218__A4 _06324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15081__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09556_ _03764_ mod.u_cpu.rf_ram.memory\[573\]\[1\] _03772_ _03777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_43_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_197_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10437__A1 _04272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08507_ _01540_ mod.u_cpu.rf_ram.memory\[326\]\[1\] _02813_ _02453_ _02814_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_145_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14649__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_196_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_212_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09487_ _03712_ _03713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_62_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07302__A1 _01608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_212_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08438_ mod.u_cpu.rf_ram.memory\[388\]\[1\] mod.u_cpu.rf_ram.memory\[389\]\[1\] mod.u_cpu.rf_ram.memory\[390\]\[1\]
+ mod.u_cpu.rf_ram.memory\[391\]\[1\] _02020_ _01995_ _02745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_106_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_197_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_225_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_156_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_211_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_183_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13926__A2 _06901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_184_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08369_ _02668_ _02671_ _02675_ _01687_ _02676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__14799__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10400_ _04392_ _00311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_11380_ _05046_ mod.u_cpu.rf_ram.memory\[302\]\[0\] _05059_ _05060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_178_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10331_ _04176_ _04344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_109_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07718__I _01757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_180_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13050_ _06199_ mod.u_cpu.rf_ram.memory\[79\]\[1\] _06201_ _06203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_10262_ _04186_ _04295_ _04296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_180_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12001_ _05483_ _05484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_133_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10193_ _03737_ _04247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_78_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07464__S1 _01771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11176__S _04919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10080__S _04165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13952_ _03430_ _03433_ _03438_ _06925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_87_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08869__A1 _02542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_235_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15424__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12903_ _06091_ _01115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_246_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09530__A2 _03717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13883_ _06468_ _06874_ _06875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_207_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_207_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15622_ _01393_ net3 mod.u_cpu.cpu.ctrl.i_jump vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12834_ _06045_ _01092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2030 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_262_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2041 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2052 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_265_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_234_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_222_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2063 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_215_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2074 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_215_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15553_ _01324_ net3 mod.u_cpu.cpu.decode.opcode\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15574__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2085 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12765_ _03950_ _05978_ _06000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2096 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14504_ _00358_ net3 mod.u_cpu.rf_ram.memory\[435\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_230_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11716_ _05249_ _05287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_187_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15484_ _01255_ net3 mod.u_arbiter.i_wb_cpu_dbus_adr\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12696_ _05955_ _01044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_226_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_230_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_187_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14435_ _00289_ net3 mod.u_cpu.rf_ram.memory\[470\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_187_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11647_ _04195_ _05239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13917__A2 _06791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09046__A1 _03349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11928__A1 _02192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14366_ _00220_ net3 mod.u_cpu.rf_ram.memory\[504\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11578_ _05193_ _00688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_128_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13317_ _03271_ _06358_ _06411_ _06414_ _01206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_182_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10451__I1 mod.u_cpu.rf_ram.memory\[450\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10529_ _04184_ _04447_ _04479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_14297_ _00151_ net3 mod.u_cpu.rf_ram.memory\[53\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_109_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09349__A2 _03590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13248_ _06349_ _01202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_44_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13793__C _06776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13179_ _06122_ mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat\[12\] _06286_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_123_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09843__I _04002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08887__C _02467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12105__A1 _03850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07780__A1 _02083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07740_ _02047_ _02048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_111_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_266_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_238_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07363__I _01537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11703__I1 mod.u_cpu.rf_ram.memory\[252\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12900__I0 _06088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_265_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07671_ _01914_ _01979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_65_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09410_ _03642_ _03638_ _03645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_25_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12408__A2 _05757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13605__A1 _03362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_213_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_197_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10419__A1 _04311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09341_ _03386_ mod.u_scanchain_local.module_data_in\[54\] _03401_ mod.u_arbiter.i_wb_cpu_dbus_adr\[17\]
+ _03587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_244_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09272_ _03488_ _03528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__14941__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07391__S0 _01697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11219__I0 _04936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08223_ _02527_ mod.u_cpu.rf_ram.memory\[516\]\[0\] _02530_ _02531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09037__A1 _03337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_193_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14030__A1 mod.u_arbiter.i_wb_cpu_rdt\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12645__S _05921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11919__A1 _05428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08154_ _02116_ _02462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_174_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08085_ _02126_ _02393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_146_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12195__I1 mod.u_cpu.rf_ram.memory\[202\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_255_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07982__B _02289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_103_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14321__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_130_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15447__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09753__I _03932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4905 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08987_ _03281_ _03283_ _03285_ _03291_ _03292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XFILLER_76_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07771__A1 _02039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4916 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4927 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4938 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07938_ mod.u_cpu.rf_ram.memory\[237\]\[0\] _02246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_4949 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13844__A1 _06367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_257_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_228_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_186_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08166__I3 mod.u_cpu.rf_ram.memory\[555\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14471__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15597__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07869_ _02157_ _02176_ _02177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_83_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09608_ _03787_ _03818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_71_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_244_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10880_ _04716_ _00467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_216_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11458__I0 _05096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__13224__B _06330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09539_ _03761_ _03762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__12619__I _05886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09276__A1 _03528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_262_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_223_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_197_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12550_ _05806_ _05858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_197_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_240_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_185_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07382__S0 _01689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_11501_ _05128_ mod.u_cpu.rf_ram.memory\[283\]\[1\] _05140_ _05142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_212_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_197_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_156_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_169_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12481_ _05657_ _04309_ _05814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_14220_ _03735_ mod.u_cpu.rf_ram.memory\[249\]\[1\] _07106_ _07108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_123_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11432_ _04817_ _05093_ _05094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_138_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09579__A2 _03786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07876__C _02166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14151_ _02261_ _07064_ _07065_ _01389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_4_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11363_ _05046_ mod.u_cpu.rf_ram.memory\[305\]\[0\] _05048_ _05049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_153_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13102_ _06236_ _06237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_10314_ _04333_ _00284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_113_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14082_ _06577_ _07021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_11294_ _04978_ mod.u_cpu.rf_ram.memory\[316\]\[0\] _05001_ _05002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_65_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08988__B _03256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13033_ _06184_ mod.u_cpu.rf_ram.memory\[108\]\[1\] _06190_ _06192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_106_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07892__B _01714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10245_ _04267_ mod.u_cpu.rf_ram.memory\[482\]\[1\] _04282_ _04284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_152_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08634__S0 _02092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_266_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_154_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_266_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10176_ _04217_ mod.u_cpu.rf_ram.memory\[492\]\[0\] _04235_ _04236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_120_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14088__A1 _03836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14814__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08500__C _01870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_248_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14984_ _00838_ net3 mod.u_cpu.rf_ram.memory\[61\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_130_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_208_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09503__A2 _03728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13935_ _06909_ _06910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_130_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_247_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_250_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13866_ _06791_ _06672_ _06858_ _06859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_62_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_263_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__14964__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15605_ _01376_ net3 mod.u_cpu.rf_ram.memory\[87\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12817_ _06034_ _01086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_188_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13797_ _06383_ _06364_ _06790_ _06395_ _06797_ _06798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_62_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15536_ _01307_ net3 mod.u_cpu.cpu.immdec.imm30_25\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_203_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12748_ _05395_ _05422_ _05989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_203_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08943__S _01478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_176_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_230_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_15467_ _01241_ net3 mod.u_cpu.cpu.ctrl.o_ibus_adr\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__14012__A1 _03458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12679_ _05312_ _05940_ _05944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_175_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09838__I _03889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14418_ _00272_ net3 mod.u_cpu.rf_ram.memory\[478\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_15398_ _01173_ net3 mod.u_cpu.rf_ram.memory\[100\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_239_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14349_ _00203_ net3 mod.u_cpu.rf_ram.memory\[513\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_183_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14344__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08898__B _02520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08910_ mod.u_cpu.rf_ram.memory\[525\]\[1\] _03217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_103_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09890_ _02567_ _04034_ _04035_ _00158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10188__I0 _04217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_170_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09573__I _03790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_257_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10888__A1 _04389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08841_ mod.u_cpu.rf_ram.memory\[45\]\[1\] _03148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__14494__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07753__A1 _02057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_250_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08772_ mod.u_cpu.rf_ram.memory\[117\]\[1\] _03079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13826__A1 _06471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_239_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07723_ _01857_ mod.u_cpu.rf_ram.memory\[270\]\[0\] _02029_ _02030_ _02031_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__08928__S1 _02543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_226_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07654_ _01752_ _01962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_198_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_240_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_41_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07585_ _01856_ _01893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_53_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13054__A2 _06193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_179_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09324_ _03436_ mod.u_scanchain_local.module_data_in\[51\] _03402_ mod.u_arbiter.i_wb_cpu_dbus_adr\[14\]
+ _03573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_222_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_167_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_194_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12801__A2 _06011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_179_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10812__A1 _04668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_194_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09255_ _03507_ _03508_ _03503_ _03514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__14003__A1 mod.u_arbiter.i_wb_cpu_rdt\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14003__B2 mod.u_arbiter.i_wb_cpu_dbus_dat\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09748__I _03928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08206_ _02484_ _02513_ _02514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09186_ mod.u_arbiter.i_wb_cpu_rdt\[19\] mod.u_arbiter.i_wb_cpu_dbus_dat\[16\] _03464_
+ _03465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__13357__A3 _06452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08608__I1 mod.u_cpu.rf_ram.memory\[129\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13601__I1 _03899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11612__I0 _05199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08137_ _02337_ _02425_ _02444_ _01591_ _02445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_181_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09430__A1 _03659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08233__A2 _02524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_175_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08084__I2 _02389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_218_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10040__A2 _04137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08068_ _02352_ _02372_ _02375_ _02361_ _02376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_150_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12317__A1 _05515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14837__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13365__I0 _03664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07992__A1 _02298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12868__A2 _04687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10030_ _04117_ mod.u_cpu.rf_ram.memory\[512\]\[0\] _04129_ _04130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_5414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07744__A1 _02046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08320__C _01742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13817__A1 _06423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14987__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_263_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08919__S1 _02495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_229_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11981_ _05422_ _05471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_72_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13720_ _06726_ _06314_ _06725_ _06441_ _06727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_72_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_217_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_205_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10932_ _04751_ _00484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_245_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_232_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07731__I _01485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_232_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13651_ _06661_ _06662_ _06663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_182_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10863_ _04700_ _04704_ _04705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_12602_ _03796_ _05882_ _05893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_158_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13582_ _06611_ _01274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_10794_ _04641_ mod.u_cpu.rf_ram.memory\[394\]\[1\] _04655_ _04657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XPHY_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_200_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_158_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_185_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_15321_ mod.u_cpu.rf_ram_if.rtrig0 net3 mod.u_cpu.rf_ram_if.rtrig1 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_12533_ _01775_ _05846_ _05847_ _00989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_212_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_184_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__11851__I0 _05364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__14367__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_200_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09658__I _03857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15252_ _00077_ net4 mod.u_arbiter.i_wb_cpu_rdt\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_32_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__15612__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12464_ _05790_ _05799_ _05801_ _03686_ _05802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_123_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14203_ _06152_ _06150_ _07098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11415_ _05071_ mod.u_cpu.rf_ram.memory\[296\]\[0\] _05082_ _05083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_172_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13753__B1 _06283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_15183_ _01036_ net3 mod.u_cpu.rf_ram.memory\[121\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_153_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12395_ _05749_ _00949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09421__A1 _03496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07178__I _01485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_193_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14134_ _07054_ _01383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_11346_ _05036_ _00613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_193_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_181_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12308__A1 _04873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14065_ mod.u_arbiter.i_wb_cpu_dbus_dat\[31\] _06919_ _07010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11277_ _04988_ _04989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09024__I1 mod.u_arbiter.i_wb_cpu_dbus_dat\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_239_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13016_ _06180_ _01139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_10228_ _03960_ _04272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_228_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_255_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13808__A1 _06418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10159_ _04221_ _00241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_66_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10590__I0 _04506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13808__B2 _06442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_181_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14967_ _00821_ net3 mod.u_cpu.rf_ram.memory\[215\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_47_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12331__I1 mod.u_cpu.rf_ram.memory\[184\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_208_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13918_ _06451_ _06874_ _06487_ _06814_ _06897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_251_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14898_ _00752_ net3 mod.u_cpu.rf_ram.memory\[235\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07641__I _01758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08160__A1 _02455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_222_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07594__S0 _01841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13849_ _06739_ mod.u_arbiter.i_wb_cpu_rdt\[5\] _06455_ _06843_ _06844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_35_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15142__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13036__A2 _06193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__12095__I0 _05533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07370_ _01677_ _01678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_210_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_204_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11598__A2 _05191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_176_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15519_ _01290_ net3 mod.u_cpu.cpu.genblk3.csr.timer_irq_r vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_30_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_198_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15292__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09040_ mod.u_cpu.cpu.state.o_cnt_r\[3\] _03342_ _03259_ _03343_ _03344_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_191_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_117_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_15_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12547__A1 _05649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_191_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13744__B1 _06338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_129_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09412__A1 _03439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09942_ _04017_ _04071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_131_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07816__I _01687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09873_ _03915_ _04023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07726__A1 _01740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11338__I _04795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_219_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11522__A2 _03791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4009 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08824_ mod.u_cpu.rf_ram.memory\[16\]\[1\] mod.u_cpu.rf_ram.memory\[17\]\[1\] mod.u_cpu.rf_ram.memory\[18\]\[1\]
+ mod.u_cpu.rf_ram.memory\[19\]\[1\] _02403_ _02367_ _03131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_258_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_245_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08755_ _02532_ mod.u_cpu.rf_ram.memory\[100\]\[1\] _03061_ _03062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_73_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13275__A2 _06360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07706_ _01998_ mod.u_cpu.rf_ram.memory\[260\]\[0\] _02013_ _02014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_2618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_214_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_241_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_227_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08686_ mod.u_cpu.rf_ram.memory\[206\]\[1\] mod.u_cpu.rf_ram.memory\[207\]\[1\] _01545_
+ _02993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10333__I0 _04345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08151__A1 _02457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1906 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_241_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_226_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_199_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_198_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1917 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_199_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07637_ mod.u_cpu.rf_ram.memory\[288\]\[0\] mod.u_cpu.rf_ram.memory\[289\]\[0\] mod.u_cpu.rf_ram.memory\[290\]\[0\]
+ mod.u_cpu.rf_ram.memory\[291\]\[0\] _01774_ _01932_ _01945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_1928 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1939 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_183_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09679__S _03874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_224_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07568_ mod.u_cpu.rf_ram.memory\[373\]\[0\] _01876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__15635__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09307_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[13\] _03557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__10636__I1 mod.u_cpu.rf_ram.memory\[420\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_179_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07499_ _01806_ _01807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_142_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_194_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09238_ _03498_ _03499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_21_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10261__A2 _04068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_210_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13929__S _06901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_181_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09169_ _03454_ _00014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09403__A1 _03614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08837__S0 _02406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11200_ _04935_ _00568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_107_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11210__A1 _04804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12180_ _05583_ mod.u_cpu.rf_ram.memory\[204\]\[1\] _05601_ _05603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_135_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13728__I _06494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_190_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11131_ _04880_ mod.u_cpu.rf_ram.memory\[342\]\[1\] _04888_ _04890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__15015__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11062_ _04796_ _04841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_135_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_5222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07717__A1 _02022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_237_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10013_ _03969_ _04118_ _04119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_114_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xtiny_user_project_103 la_data_out[21] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_118_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xtiny_user_project_114 la_data_out[32] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_5255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_125 la_data_out[43] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_5277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xtiny_user_project_136 la_data_out[54] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__08390__A1 _02272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtiny_user_project_147 user_irq[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_5288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14821_ _00675_ net3 mod.u_cpu.rf_ram.memory\[277\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_95_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_158 wbs_dat_o[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_5299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15165__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_4565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xtiny_user_project_169 wbs_dat_o[19] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_64_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11184__S _04923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14752_ _00606_ net3 mod.u_cpu.rf_ram.memory\[311\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_151_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_217_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_151_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11964_ _05442_ mod.u_cpu.rf_ram.memory\[539\]\[0\] _05459_ _05460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10324__I0 _04326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_233_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_205_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_204_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_205_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09190__I0 mod.u_arbiter.i_wb_cpu_rdt\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13703_ _06371_ _06389_ _06711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_3897 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12079__I _03841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10915_ _04739_ mod.u_cpu.rf_ram.memory\[375\]\[1\] _04737_ _04740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_14683_ _00537_ net3 mod.u_cpu.rf_ram.memory\[346\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11895_ _05411_ _00787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13018__A2 _03919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_220_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12077__I0 _05533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13634_ _06455_ _06647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_60_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10846_ _04679_ mod.u_cpu.rf_ram.memory\[385\]\[0\] _04691_ _04692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_60_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_220_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_198_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_201_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11824__I0 _05350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13565_ mod.u_arbiter.i_wb_cpu_dbus_adr\[16\] mod.u_arbiter.i_wb_cpu_dbus_adr\[17\]
+ _06599_ _06602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_12_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10777_ _04646_ _00434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_197_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11711__I _03803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15304_ _00065_ net4 mod.u_scanchain_local.module_data_in\[61\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_157_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12516_ _02137_ _05835_ _05836_ _00983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_199_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13496_ _03635_ _06551_ _06552_ _03642_ _06556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_139_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15235_ _01088_ net3 mod.u_cpu.rf_ram.memory\[126\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_157_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12447_ _03412_ _03400_ _05785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_173_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15166_ _01019_ net3 mod.u_cpu.rf_ram.memory\[151\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12378_ _05738_ _00943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_125_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07956__A1 _02174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14117_ _06181_ _03911_ _07044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_4_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11329_ _04741_ _05011_ _05025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_114_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15097_ _00951_ net3 mod.u_cpu.rf_ram.memory\[479\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_141_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14048_ _06963_ _06998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_141_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15508__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13574__S _06604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10563__I0 _04498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_227_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08895__C _02487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__10997__I _04795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_208_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08540_ _01807_ mod.u_cpu.rf_ram.memory\[292\]\[1\] _02846_ _02847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_78_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__14532__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_209_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10315__I0 _04330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08133__A1 _02161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07371__I _01660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09181__I0 mod.u_arbiter.i_wb_cpu_rdt\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_223_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08471_ _01991_ _02778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_51_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14206__A1 _06047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_243_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11822__S _05359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07422_ mod.u_cpu.rf_ram.memory\[407\]\[0\] _01730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_196_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_211_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_206_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14682__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07353_ _01660_ _01661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_176_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09633__A1 _03775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11621__I _04959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_206_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_52_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15240__D _01093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_206_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_143_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07284_ _01445_ _01592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_108_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08135__C _02185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09023_ _03306_ _03269_ _03268_ _03328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_191_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15038__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_191_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09397__B1 _03401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07546__I _01499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09925_ _04013_ _03843_ _04059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_131_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__15188__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09856_ _04011_ _00148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_252_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08807_ _03102_ _03104_ _03113_ _02664_ _03114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_105_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09787_ _03870_ _03939_ _03959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_2_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_234_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13283__I _06380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_215_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08738_ _02632_ mod.u_cpu.rf_ram.memory\[254\]\[1\] _03044_ _01702_ _03045_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_3149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_215_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08124__A1 _02410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08669_ _02711_ _02974_ _02975_ _01723_ _02976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XTAP_1725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12828__S _06040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11732__S _05297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_202_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10700_ _04594_ _00409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_230_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_202_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12059__I0 _05521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_202_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11680_ _05253_ _05262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10482__A2 _04447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__12759__A1 _04668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_201_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10631_ _04414_ _04548_ _04549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_195_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11531__I _05107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11431__A1 _04412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13350_ _06358_ _06419_ _06420_ _06446_ _01207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_210_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11282__I1 mod.u_cpu.rf_ram.memory\[318\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10562_ _04501_ _00364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_155_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13708__B1 _06713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12301_ _05685_ _00919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11982__A2 _05471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_212_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_182_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13281_ _03501_ mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat\[1\] _06378_ _06379_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_6_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10493_ _04450_ mod.u_cpu.rf_ram.memory\[444\]\[1\] _04454_ _04456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_154_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15020_ _00874_ net3 mod.u_cpu.rf_ram.memory\[73\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_170_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13184__A1 _05783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12232_ mod.u_cpu.rf_ram.memory\[197\]\[1\] _05617_ _05637_ _05639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_108_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__14405__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12163_ mod.u_cpu.rf_ram.memory\[73\]\[1\] _05468_ _05590_ _05592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_146_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11114_ _04864_ mod.u_cpu.rf_ram.memory\[344\]\[0\] _04877_ _04878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_151_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12094_ _05545_ _00852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_151_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_20 io_oeb[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__08996__B _03300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11907__S _05418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12534__I1 _05765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_31 io_oeb[23] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_5030 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11498__A1 _05139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11045_ _04825_ mod.u_cpu.rf_ram.memory\[355\]\[1\] _04828_ _04830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_89_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5041 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_231_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_42 io_oeb[34] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_1_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14555__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5052 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_162_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_53 io_out[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__10545__I0 _04481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_209_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xtiny_user_project_64 io_out[20] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__08363__A1 _01561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_264_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5063 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xtiny_user_project_75 io_out[31] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_5074 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xtiny_user_project_86 la_data_out[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_5085 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5096 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xtiny_user_project_97 la_data_out[15] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_4362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_237_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_218_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14804_ _00658_ net3 mod.u_cpu.rf_ram.memory\[285\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_91_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12298__I0 _05679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_252_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08287__I _02030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12996_ mod.u_cpu.cpu.genblk3.csr.mcause3_0\[2\] _06167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_218_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_205_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14735_ _00589_ net3 mod.u_cpu.rf_ram.memory\[320\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11947_ _05448_ _05447_ _05449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_91_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_205_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_229_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2960 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_205_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_178_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2971 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_221_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_206_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_178_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2982 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11670__A1 _04868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14666_ _00520_ net3 mod.u_cpu.rf_ram.memory\[354\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2993 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11878_ _02357_ _05398_ _05399_ _00782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_178_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_207_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13617_ _01926_ _06633_ _06634_ _01286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_60_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10258__S _04291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10829_ _04679_ mod.u_cpu.rf_ram.memory\[388\]\[0\] _04680_ _04681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09615__A1 _03775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14597_ _00451_ net3 mod.u_cpu.rf_ram.memory\[38\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_158_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10225__A2 _04269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13548_ _06592_ _01259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_185_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08969__A3 mod.u_cpu.cpu.csr_d_sel vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_201_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12981__B _06056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13479_ _06539_ _06546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_127_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15218_ _01071_ net3 mod.u_cpu.rf_ram.memory\[133\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_154_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__11089__S _04860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15330__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_236_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15149_ _01002_ net3 mod.u_cpu.rf_ram.memory\[160\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_142_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10784__I0 _04641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_259_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07971_ _01739_ _02256_ _02278_ _02279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_113_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09710_ _03899_ _03897_ _03900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_256_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10536__I0 _04469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07157__A2 _01465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08354__A1 _02654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15480__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09581__I _03796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09641_ _03802_ mod.u_cpu.rf_ram.memory\[564\]\[0\] _03844_ _03845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_255_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_222_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_209_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12289__I0 _05677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09572_ _03789_ _03790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08106__A1 _02410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09154__I0 mod.u_arbiter.i_wb_cpu_rdt\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_247_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_236_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08523_ _01864_ _02829_ _02830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_36_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12648__S _05921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_224_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09854__A1 _03782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08657__A2 _02963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08454_ mod.u_cpu.rf_ram.memory\[381\]\[1\] _02761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_168_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07969__C _02207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07960__S0 _02266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13789__I0 mod.u_arbiter.i_wb_cpu_rdt\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07405_ _01711_ _01712_ _01713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_56_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_196_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08385_ _02220_ _02692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_177_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07336_ _01494_ _01644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10216__A2 _04263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_221_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_221_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14428__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07267_ _01573_ _01574_ _01575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_164_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09006_ _03306_ _03307_ _03310_ _03311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__11016__I1 mod.u_cpu.rf_ram.memory\[35\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07198_ mod.u_cpu.raddr\[0\] _01506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_145_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_254_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_191_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12182__I _05309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14578__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07276__I _01528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_219_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08593__A1 _01979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11727__S _05294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09908_ _04023_ mod.u_cpu.rf_ram.memory\[532\]\[0\] _04047_ _04048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10527__I0 _04467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14103__S _07033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07779__S0 _02085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08345__A1 _02631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__12141__A2 _05576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09839_ _03999_ mod.u_cpu.rf_ram.memory\[543\]\[1\] _03997_ _04000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_111_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_207_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12850_ _02505_ _06054_ _06055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_234_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11801_ _05329_ mod.u_cpu.rf_ram.memory\[232\]\[1\] _05344_ _05346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_2234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_261_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_162_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12781_ _05962_ _06010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_1511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_215_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_54_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14520_ _00374_ net3 mod.u_cpu.rf_ram.memory\[427\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11732_ _05289_ mod.u_cpu.rf_ram.memory\[241\]\[0\] _05297_ _05298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_203_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_226_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_199_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15203__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_2289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_230_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_202_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_187_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14451_ _00305_ net3 mod.u_cpu.rf_ram.memory\[462\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11663_ _05249_ _05250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_14_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13402_ _06381_ _06439_ _06495_ _06496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_122_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10614_ _04497_ _04537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_168_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_14382_ _00236_ net3 mod.u_cpu.rf_ram.memory\[496\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__13897__B _06856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11594_ _05199_ mod.u_cpu.rf_ram.memory\[267\]\[0\] _05203_ _05204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_183_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07703__S0 _01994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13333_ _06318_ _06428_ _06429_ _06430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__15353__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10545_ _04481_ mod.u_cpu.rf_ram.memory\[435\]\[1\] _04488_ _04490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_183_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_196_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_182_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12204__I0 _05605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13264_ _06361_ _06362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_108_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10476_ _04299_ _04443_ _04444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_182_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15003_ _00857_ net3 mod.u_cpu.rf_ram.memory\[211\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_136_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12215_ _05605_ mod.u_cpu.rf_ram.memory\[198\]\[0\] _05626_ _05627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_237_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14224__D _00000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13195_ _06126_ mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat\[13\] _06302_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08584__A1 _01997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07186__I mod.u_cpu.raddr\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12146_ _05187_ _05552_ _05580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_150_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12077_ _05533_ mod.u_cpu.rf_ram.memory\[64\]\[1\] _05531_ _05534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_110_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08336__A1 _02631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_265_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11028_ _04817_ _04816_ _04818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_110_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_237_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11436__I _05045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08887__A2 _03190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__13880__A2 _06871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_266_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__11891__A1 _05408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_253_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xtiny_user_project_8 io_oeb[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_18_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09836__A1 _03945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12979_ _01453_ _06152_ _06153_ _06154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XTAP_3491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13632__A2 _06324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_244_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_45_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_206_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14718_ _00572_ net3 mod.u_cpu.rf_ram.memory\[328\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_61_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07311__A2 _01606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_220_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14649_ _00503_ net3 mod.u_cpu.rf_ram.memory\[363\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_162_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11171__I _04879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_203_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13396__A1 _06483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08170_ _02477_ _02478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_53_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09064__A2 _03363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_174_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07121_ mod.u_cpu.cpu.csr_d_sel _01430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_203_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14720__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13699__A2 _06704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08413__C _01678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08575__A1 _01981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10382__A1 _04225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14870__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07954_ _02180_ _02261_ _02262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_173_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_228_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07885_ _01682_ mod.u_cpu.rf_ram.memory\[220\]\[0\] _02193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08878__A2 _03177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_229_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09624_ _03831_ _00096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_83_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11882__A1 _04965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15226__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10685__A2 _04575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14120__I0 _07041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09555_ _02497_ _03772_ _03776_ _00082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_83_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_243_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08506_ _02672_ _02812_ _02813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_93_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_212_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_145_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09486_ _03702_ _03711_ _03712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__12682__I0 _05938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_224_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_212_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_196_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_168_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14250__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15376__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08437_ _01680_ _02743_ _02744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_196_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_196_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09687__S _03880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_196_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08368_ _01567_ mod.u_cpu.rf_ram.memory\[486\]\[1\] _02674_ _02109_ _02675_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_183_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07319_ _01577_ mod.u_cpu.rf_ram.memory\[486\]\[0\] _01626_ _01582_ _01627_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_20_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_192_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08299_ _01533_ _02606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_178_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_165_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10330_ _04343_ _00290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_192_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_152_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10261_ _04294_ _04068_ _04295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_117_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10748__I0 _04626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12000_ _05404_ _05483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08566__A1 _01791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10192_ _04246_ _00249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_120_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_191_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_266_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_232_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08318__A1 _02115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07734__I _01499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_247_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_13951_ _06923_ _06924_ _01330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_115_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_219_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08869__A2 _03168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13862__A2 _06849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10160__I mod.u_cpu.cpu.immdec.imm11_7\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_235_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_86_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12902_ _06086_ mod.u_cpu.rf_ram.memory\[96\]\[1\] _06089_ _06091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_13882_ _06858_ _06873_ _06874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_185_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__14111__I0 _07021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12833_ _06038_ mod.u_cpu.rf_ram.memory\[124\]\[1\] _06043_ _06045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_2020 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15621_ _01392_ net3 mod.u_cpu.cpu.bufreg2.i_cnt_done vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2031 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2042 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13614__A2 _03378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2053 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2064 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15552_ _01323_ net3 mod.u_cpu.cpu.decode.opcode\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12764_ _05999_ _01068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2075 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2086 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2097 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11715_ _05286_ _00732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_203_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_199_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14503_ _00357_ net3 mod.u_cpu.rf_ram.memory\[436\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_30_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_203_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15483_ _01254_ net3 mod.u_arbiter.i_wb_cpu_dbus_adr\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_202_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12695_ mod.u_cpu.rf_ram.memory\[141\]\[1\] _05950_ _05953_ _05955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_230_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_203_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11646_ _05238_ _00711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__14743__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14434_ _00288_ net3 mod.u_cpu.rf_ram.memory\[470\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12425__I0 _05761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_204_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11928__A2 _05434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12050__A1 _05515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14365_ _00219_ net3 mod.u_cpu.rf_ram.memory\[505\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11577_ _05180_ mod.u_cpu.rf_ram.memory\[270\]\[0\] _05192_ _05193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_156_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_196_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14178__I0 _07057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13316_ mod.u_cpu.cpu.immdec.imm11_7\[1\] _06413_ _06357_ _06414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_10_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10528_ _04478_ _00353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_170_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14296_ _00150_ net3 mod.u_cpu.rf_ram.memory\[53\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_122_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14893__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08233__C _02469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10335__I _04247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13247_ _06273_ mod.u_cpu.rf_ram.memory\[92\]\[0\] _06348_ _06349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12751__S _05989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10459_ _04431_ _00331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_100_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13178_ _06284_ _06285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_124_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_123_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13646__I _06655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12129_ _05300_ _05568_ _05569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_112_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15249__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08309__A1 _02532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12105__A2 _05552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_250_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_226_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13853__A2 _06836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07670_ _01832_ _01978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10667__A2 _04571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_203_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14273__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_225_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__15399__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12198__S _05615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_252_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09340_ _03571_ _03585_ _03586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__11616__A1 _04539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09285__A2 _03538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09271_ _03506_ _03526_ _03527_ _00046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_221_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_205_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11830__S _05362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08222_ _02528_ _02529_ _02530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07391__S1 _01698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_148_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11919__A2 _05423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08153_ _02115_ _02461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_140_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_146_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07819__I _02126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08084_ _02384_ _02387_ _02389_ _02390_ _02391_ _01720_ _02392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_147_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07982__C _02141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10355__A1 _04360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_102_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_251_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_130_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08986_ _03289_ _03290_ _03291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_102_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_229_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4906 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07554__I _01509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4917 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4928 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_229_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07937_ _01681_ _02245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10107__A1 _04184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4939 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14616__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11076__I _03750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_256_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07868_ mod.u_cpu.rf_ram.memory\[205\]\[0\] _02176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_29_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08720__A1 _01698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09607_ _03817_ _00093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_3_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_249_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_204_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07799_ _01854_ _02107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11804__I _05132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09538_ _03732_ _03761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__14766__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11458__I1 mod.u_cpu.rf_ram.memory\[28\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08385__I _02220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_145_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_227_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_212_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07287__A1 _01573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09469_ mod.u_cpu.rf_ram_if.wdata1_r\[0\] mod.u_cpu.rf_ram_if.wdata0_r _01449_ _03695_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07222__C _01529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12280__A1 _05428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_212_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_200_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_11500_ _05141_ _00662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_157_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07382__S1 _01683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_185_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12480_ _05812_ _05813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_200_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_200_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09210__S _03474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11431_ _04412_ _05062_ _05093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__10356__S _04361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_123_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10969__I0 _04774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_193_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08787__A1 _01662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14150_ _07026_ _07064_ _07065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__13780__A1 _06494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11362_ _05047_ _05038_ _05048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_125_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13101_ _06017_ _06236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_164_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10313_ _04326_ mod.u_cpu.rf_ram.memory\[472\]\[0\] _04332_ _04333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_98_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14081_ _07020_ _01364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_11293_ _04859_ _04990_ _05001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_180_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08539__A1 _01843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13032_ _06191_ _01144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_10244_ _04283_ _00264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_4_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13466__I _06509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08634__S1 _02098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_234_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_105_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_191_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10175_ _04233_ _04234_ _04235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_67_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14088__A2 _05279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09880__S _04027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14296__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14983_ _00837_ net3 mod.u_cpu.rf_ram.memory\[213\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_47_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_266_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15541__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13835__A2 _03682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_208_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13934_ _03394_ _03280_ _06907_ _06908_ _05800_ _06909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_35_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_207_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_13865_ _06282_ _06294_ _06305_ _06858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_262_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_234_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_216_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15604_ _01375_ net3 mod.u_cpu.rf_ram.memory\[87\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__13599__A1 _03694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12816_ _06019_ mod.u_cpu.rf_ram.memory\[127\]\[1\] _06031_ _06034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__13599__B2 _03659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13796_ _06321_ _06683_ _06797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_163_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_250_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_231_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15535_ _01306_ net3 mod.u_cpu.cpu.immdec.imm30_25\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_37_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12747_ _05988_ _01062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12746__S _05986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_231_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_179_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12678_ _05943_ _01038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_15466_ _01240_ net3 mod.u_cpu.cpu.ctrl.o_ibus_adr\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_187_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__14012__A2 _06964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12023__A1 _05452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11629_ _05226_ _05210_ _05227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_14417_ _00271_ net3 mod.u_cpu.rf_ram.memory\[47\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_204_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_200_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15397_ _01172_ net3 mod.u_cpu.rf_ram.memory\[100\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_129_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_184_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08617__I2 mod.u_cpu.rf_ram.memory\[138\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08778__A1 _02325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_190_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_184_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13771__A1 _06415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_200_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14348_ _00202_ net3 mod.u_cpu.rf_ram.memory\[513\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_116_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14279_ _00133_ net3 mod.u_cpu.rf_ram.memory\[548\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_83_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15071__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10337__A1 _04189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_170_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10188__I1 mod.u_cpu.rf_ram.memory\[490\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14639__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_170_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08840_ mod.u_cpu.rf_ram.memory\[46\]\[1\] mod.u_cpu.rf_ram.memory\[47\]\[1\] _01577_
+ _03147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10888__A2 _04108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_258_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07753__A2 _02060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08771_ mod.u_cpu.rf_ram.memory\[112\]\[1\] mod.u_cpu.rf_ram.memory\[113\]\[1\] mod.u_cpu.rf_ram.memory\[114\]\[1\]
+ mod.u_cpu.rf_ram.memory\[115\]\[1\] _01664_ _02323_ _03078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_215_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13826__A2 _06823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_257_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_238_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07722_ _01782_ _02030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_266_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__14789__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_254_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08702__A1 _02665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07505__A2 _01801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07653_ _01960_ _01961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_226_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_214_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_253_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07584_ mod.u_cpu.rf_ram.memory\[360\]\[0\] mod.u_cpu.rf_ram.memory\[361\]\[0\] mod.u_cpu.rf_ram.memory\[362\]\[0\]
+ mod.u_cpu.rf_ram.memory\[363\]\[0\] _01843_ _01838_ _01892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__12637__I0 _05904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09323_ _03569_ _03571_ _03572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_178_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_240_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11560__S _05181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09254_ _03506_ _03512_ _03513_ _00043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_179_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10812__A2 _04669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_193_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14003__A2 _06964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08205_ mod.u_cpu.rf_ram.memory\[567\]\[0\] _02513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_166_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09185_ _03451_ _03464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_239_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08769__A1 _02283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08313__S0 _02593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08136_ _02149_ _02434_ _02443_ _02444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__15414__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13762__A1 _03298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_175_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_190_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09430__A2 _03402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08084__I3 _02390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08067_ _02356_ mod.u_cpu.rf_ram.memory\[78\]\[0\] _02374_ _02359_ _02375_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_49_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09764__I _03941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13365__I1 _03663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13514__A1 mod.u_cpu.cpu.state.o_cnt_r\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_255_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10328__A1 _04251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11376__I0 _05050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15564__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08601__C _01631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_102_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07744__A2 _02050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_216_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13278__B1 _06370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08969_ _01421_ mod.u_cpu.cpu.branch_op mod.u_cpu.cpu.csr_d_sel _03274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_130_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_257_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11980_ _05412_ _05470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__14111__S _07039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_217_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10931_ _04728_ mod.u_cpu.rf_ram.memory\[372\]\[0\] _04750_ _04751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_90_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_244_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_205_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_216_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13650_ _06320_ _06368_ _06662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_140_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10862_ _04703_ _04704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_147_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_262_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12601_ _05892_ _01012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_242_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13581_ mod.u_arbiter.i_wb_cpu_dbus_adr\[23\] mod.u_arbiter.i_wb_cpu_dbus_adr\[24\]
+ _06609_ _06611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XPHY_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10793_ _04656_ _00440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12566__S _05866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_34_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15320_ _01099_ net3 mod.u_cpu.raddr\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12532_ _05642_ _05846_ _05847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07887__C _01833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_185_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_185_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07680__A1 _01981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15251_ _00076_ net4 mod.u_arbiter.i_wb_cpu_rdt\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12463_ _05800_ _05801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10086__S _04169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15094__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_200_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11414_ _04804_ _05058_ _05082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13753__A1 _06726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14202_ _06152_ _06151_ _07097_ _01409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__13753__B2 _06712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15182_ _01035_ net3 mod.u_cpu.rf_ram.memory\[121\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12394_ _05745_ mod.u_cpu.rf_ram.memory\[509\]\[1\] _05747_ _05749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_165_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10567__A1 _01780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14133_ _07043_ mod.u_cpu.rf_ram.memory\[115\]\[0\] _07053_ _07054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_11345_ _05032_ mod.u_cpu.rf_ram.memory\[308\]\[1\] _05034_ _05036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_193_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_180_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_154_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14064_ _07008_ _07009_ _01358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_153_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11276_ _03755_ _04701_ _04988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__10319__A1 _04311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09024__I2 mod.u_arbiter.i_wb_cpu_dbus_dat\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13015_ _06105_ mod.u_cpu.rf_ram.memory\[85\]\[1\] _06178_ _06180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_10227_ _04271_ _00259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_95_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_234_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14931__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13108__I1 _06221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10158_ _04215_ mod.u_cpu.rf_ram.memory\[494\]\[1\] _04219_ _04221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_67_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_239_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11645__S _05236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_208_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14966_ _00820_ net3 mod.u_cpu.rf_ram.memory\[215\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10089_ _04171_ _00221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_236_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07922__I _01719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13917_ _06647_ _06791_ _06640_ _06896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_223_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14897_ _00751_ net3 mod.u_cpu.rf_ram.memory\[236\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_169_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_263_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_235_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07594__S1 _01844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13848_ _06334_ mod.u_arbiter.i_wb_cpu_rdt\[21\] _06843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_50_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_251_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_204_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_245_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_200_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13779_ _06777_ _06780_ _06331_ _06781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_222_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__14311__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15518_ _01289_ net3 mod.u_cpu.rf_ram.memory\[309\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__15437__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_175_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09660__A2 _03859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_175_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15449_ _01223_ net3 mod.u_cpu.cpu.ctrl.o_ibus_adr\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_176_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07369__I _01550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_198_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13744__A1 mod.u_cpu.cpu.immdec.imm19_12_20\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12547__A2 _05831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_175_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13744__B2 _06741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_176_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__15587__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14461__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07423__A1 _01729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09941_ _02552_ _04069_ _04070_ _00174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_131_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_252_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_213_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09872_ _04022_ _00153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_219_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10030__I0 _04117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08823_ _02365_ _03122_ _03129_ _02185_ _03130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_135_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10730__A1 _04189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08754_ _02171_ _03060_ _03061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_100_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_261_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07705_ _01711_ _02012_ _02013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_94_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08685_ _02972_ _02978_ _02985_ _02991_ _01489_ _02992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XTAP_2619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_226_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1907 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07636_ _01791_ _01931_ _01943_ _01944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_1918 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08782__S0 _02249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1929 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_263_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07567_ _01825_ _01875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12235__A1 _05593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_241_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09306_ _03546_ _03553_ _03556_ _00053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__09100__A1 _03385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13983__A1 mod.u_arbiter.i_wb_cpu_rdt\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13983__B2 mod.u_arbiter.i_wb_cpu_dbus_dat\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07498_ _01603_ _01806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_146_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10797__A1 _04527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_210_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09237_ mod.u_cpu.cpu.genblk1.align.ctrl_misal _03498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__14804__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_210_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_33_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07279__I _01586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13735__A1 _06739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12538__A2 _05849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_194_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09168_ mod.u_arbiter.i_wb_cpu_rdt\[12\] mod.u_arbiter.i_wb_cpu_dbus_dat\[9\] _03452_
+ _03454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_119_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08837__S1 _02218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_181_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08119_ mod.u_cpu.rf_ram.memory\[37\]\[0\] _02427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_163_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09099_ _03399_ _03400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_108_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11130_ _04889_ _00544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_163_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14954__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_150_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11061_ _04840_ _00524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_122_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_192_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_5223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07717__A2 mod.u_cpu.rf_ram.memory\[268\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10012_ _03995_ _04118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08914__A1 _02551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_77_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xtiny_user_project_104 la_data_out[22] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_49_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_192_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_49_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xtiny_user_project_115 la_data_out[33] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_103_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_237_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_130_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_126 la_data_out[44] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_95_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_137 la_data_out[55] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_5278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14820_ _00674_ net3 mod.u_cpu.rf_ram.memory\[277\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_5289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xtiny_user_project_148 user_irq[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_64_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_159 wbs_dat_o[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_218_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_218_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_229_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14751_ _00605_ net3 mod.u_cpu.rf_ram.memory\[312\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12474__A1 _05395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_251_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11963_ _05139_ _03996_ _05459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_245_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10324__I1 mod.u_cpu.rf_ram.memory\[470\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13702_ _06710_ _01295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__14334__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_217_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10914_ _04719_ _04739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_11894_ _05406_ mod.u_cpu.rf_ram.memory\[226\]\[1\] _05409_ _05411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_3898 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14682_ _00536_ net3 mod.u_cpu.rf_ram.memory\[346\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09890__A2 _04034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_60_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_233_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07898__B _02205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13633_ mod.u_arbiter.i_wb_cpu_rdt\[31\] _03458_ _03503_ _06646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_10845_ _04285_ _04687_ _04691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_38_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_204_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10088__I0 _04157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_13564_ _06601_ _01266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_10776_ mod.u_cpu.rf_ram.memory\[397\]\[0\] _04396_ _04645_ _04646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_185_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14484__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15303_ _00064_ net4 mod.u_scanchain_local.module_data_in\[60\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12515_ _05759_ _05835_ _05836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_125_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13026__I0 _06186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_185_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07410__C _01717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13495_ _06555_ _01243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_121_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_240_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_200_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13726__A1 _06438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_195_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_12446_ _05783_ _05784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_15234_ _01087_ net3 mod.u_cpu.rf_ram.memory\[126\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_139_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07405__A1 _01711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12377_ _05729_ mod.u_cpu.rf_ram.memory\[17\]\[1\] _05736_ _05738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_158_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15165_ _01018_ net3 mod.u_cpu.rf_ram.memory\[152\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_176_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11328_ _05024_ _00607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_14116_ _06577_ _07043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_140_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15096_ _00950_ net3 mod.u_cpu.rf_ram.memory\[479\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_119_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10960__A1 _04369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13855__S _06335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10343__I _04302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11259_ _04951_ _04976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_14047_ mod.u_arbiter.i_wb_cpu_dbus_dat\[26\] _06989_ _06997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_80_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08905__A1 _02500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_228_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_209_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07652__I _01749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_243_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_208_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14949_ _00803_ net3 mod.u_cpu.rf_ram.memory\[21\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_36_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_224_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11174__I _04882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09181__I1 mod.u_arbiter.i_wb_cpu_dbus_dat\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08133__A2 mod.u_cpu.rf_ram.memory\[46\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08470_ _02765_ _02767_ _02776_ _01849_ _02777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_35_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_208_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_211_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07421_ _01519_ _01729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_90_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14827__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07892__A1 _01517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_210_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_223_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08516__S0 _02751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07352_ _01659_ _01660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13965__A1 mod.u_arbiter.i_wb_cpu_dbus_dat\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_188_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_176_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07283_ _01458_ _01591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_148_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_191_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09022_ mod.u_cpu.cpu.mem_if.signbit _03327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__14977__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_191_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09397__A1 _03386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_191_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10454__S _04427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09397__B2 mod.u_arbiter.i_wb_cpu_dbus_adr\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07947__A2 _02243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09924_ _04058_ _00169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_59_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09855_ _04001_ mod.u_cpu.rf_ram.memory\[540\]\[0\] _04010_ _04011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_219_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_258_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_213_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08806_ _02665_ _03105_ _03112_ _02677_ _03113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__14357__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09786_ _03915_ _03958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_73_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07562__I _01550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15602__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_233_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08737_ _02084_ _03043_ _03044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_227_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08124__A2 mod.u_cpu.rf_ram.memory\[38\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09321__A1 mod.u_cpu.cpu.ctrl.o_ibus_adr\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_215_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_198_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08668_ _01567_ mod.u_cpu.rf_ram.memory\[216\]\[1\] _02975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_1704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_183_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_199_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_187_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07619_ _01507_ _01926_ _01927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13256__I0 _06354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_183_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08599_ _01672_ _02905_ _02906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08607__B _02913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_186_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13956__A1 mod.u_arbiter.i_wb_cpu_rdt\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10630_ _04412_ _04528_ _04548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__13956__B2 _03438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10561_ _04486_ mod.u_cpu.rf_ram.memory\[432\]\[0\] _04500_ _04501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__13008__I0 _06107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11431__A2 _05062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_259_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12300_ _05677_ mod.u_cpu.rf_ram.memory\[187\]\[1\] _05683_ _05685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__13708__A1 _06318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13280_ _06377_ _03424_ _06378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_167_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10492_ _04455_ _00340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_108_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12231_ _02158_ _05637_ _05638_ _00896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_108_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13184__A2 mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12643__I _05919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_205_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_170_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12162_ _05591_ _00874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_135_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11259__I _04951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15132__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11990__I0 _05464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11113_ _04732_ _04869_ _04877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_12093_ _05539_ mod.u_cpu.rf_ram.memory\[66\]\[0\] _05544_ _05545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_151_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_10 io_oeb[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_5020 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11044_ _04829_ _00518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08996__C _01422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtiny_user_project_21 io_oeb[13] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_77_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_32 io_oeb[24] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_122_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_43 io_oeb[35] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_5031 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5042 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11742__I0 _05304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5053 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xtiny_user_project_54 io_out[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_5064 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_162_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_65 io_out[21] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_65_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_76 io_out[32] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_5075 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_77_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xtiny_user_project_87 la_data_out[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__15282__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5086 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xtiny_user_project_98 la_data_out[16] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__10170__A2 _04229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5097 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_225_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14803_ _00657_ net3 mod.u_cpu.rf_ram.memory\[286\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_4363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_206_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12447__A1 _03412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12995_ _03686_ _06166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_4396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14734_ _00588_ net3 mod.u_cpu.rf_ram.memory\[320\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11946_ _05132_ _05448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_206_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2950 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2961 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2972 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07874__A1 _02180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14665_ _00519_ net3 mod.u_cpu.rf_ram.memory\[355\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2983 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13247__I0 _06273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11877_ _05348_ _05398_ _05399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_2994 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_221_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_205_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08517__B _01788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13616_ _06249_ _06633_ _06634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_158_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10828_ _04272_ _04669_ _04680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_207_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14596_ _00450_ net3 mod.u_cpu.rf_ram.memory\[38\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_201_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13547_ mod.u_arbiter.i_wb_cpu_dbus_adr\[8\] mod.u_arbiter.i_wb_cpu_dbus_adr\[9\]
+ _06589_ _06592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_119_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10759_ _04633_ _00429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_187_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13478_ _06537_ _06545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13649__I _06404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_15217_ _01070_ net3 mod.u_cpu.rf_ram.memory\[134\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_86_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12429_ _01796_ _05771_ _05772_ _00960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_142_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15148_ _01001_ net3 mod.u_cpu.rf_ram.memory\[160\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_142_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07970_ _01791_ _02265_ _02277_ _02278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_173_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08679__S _01807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15079_ _00933_ net3 mod.u_cpu.rf_ram.memory\[182\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_99_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_214_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15625__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09926__I0 _04051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12686__A1 _05948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10536__I1 mod.u_cpu.rf_ram.memory\[436\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08354__A2 _02655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09640_ _03814_ _03843_ _03844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_68_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_256_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09571_ _03786_ _03788_ _03789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_215_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_209_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08522_ mod.u_cpu.rf_ram.memory\[343\]\[1\] _02829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__09154__I1 _03444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_212_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08453_ mod.u_cpu.rf_ram.memory\[382\]\[1\] mod.u_cpu.rf_ram.memory\[383\]\[1\] _02125_
+ _02760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_51_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13238__I0 _06276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_212_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_196_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11632__I _03733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_211_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07404_ mod.u_cpu.rf_ram.memory\[415\]\[0\] _01712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_211_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15005__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13938__A1 _05800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07960__S1 _02267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13789__I1 _03449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08384_ mod.u_cpu.rf_ram.memory\[416\]\[1\] mod.u_cpu.rf_ram.memory\[417\]\[1\] mod.u_cpu.rf_ram.memory\[418\]\[1\]
+ mod.u_cpu.rf_ram.memory\[419\]\[1\] _02559_ _02155_ _02691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_149_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_260_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07335_ _01604_ _01643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_176_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10472__I0 _04430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07266_ mod.u_cpu.rf_ram.memory\[469\]\[0\] _01574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09005_ _03308_ _03309_ _03310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__15155__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_192_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_191_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12463__I _05800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10184__S _04239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_247_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07197_ _01504_ _01505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13410__I0 _06354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11972__I0 _05464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08593__A2 _02899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09772__I _03766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09907_ _03843_ _04038_ _04047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_76_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10527__I1 mod.u_cpu.rf_ram.memory\[438\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11807__I _05328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08345__A2 _02644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07779__S1 _02086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09838_ _03889_ _03999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_219_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_150_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_262_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12429__A1 _01796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09769_ _02463_ _03943_ _03946_ _00126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_2202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11800_ _05345_ _00758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_132_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12780_ _06009_ _01074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09213__S _03479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_2257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_203_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11731_ _05047_ _05284_ _05297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13229__I0 mod.u_arbiter.i_wb_cpu_rdt\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_15_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_215_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__10359__S _04361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_230_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_30_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14450_ _00304_ net3 mod.u_cpu.rf_ram.memory\[462\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11662_ _05106_ _05249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_161_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08056__C _02363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13401_ _06438_ _06493_ _06494_ _06495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_10613_ _04536_ _00380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_11593_ _04930_ _05191_ _05203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_14381_ _00235_ net3 mod.u_cpu.rf_ram.memory\[497\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_211_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10463__I0 _04430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07703__S1 _02010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13332_ _06417_ _06326_ _06330_ _06429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_127_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10544_ _04489_ _00358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08900__S0 _02494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08281__A1 _02198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_196_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_182_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_41_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13469__I _06539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13263_ _06359_ _06360_ _06361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10475_ _04442_ _04443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_157_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11168__A1 _04913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_15002_ _00856_ net3 mod.u_cpu.rf_ram.memory\[211\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09883__S _04030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14522__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12214_ _05355_ _05611_ _05626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08033__A1 _01696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13194_ _06298_ _06300_ _06301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_135_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14106__A1 _07026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_233_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_12145_ _05579_ _00869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_194_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09781__A1 _03878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_111_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09908__I0 _04023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_256_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_12076_ _05483_ _05533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_155_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14672__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_2_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08336__A2 _02634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11027_ _03898_ _04817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_65_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_238_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_225_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_252_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_4193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15028__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtiny_user_project_9 io_oeb[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_206_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13093__A1 _05888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12978_ _03268_ _06153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13632__A3 _06643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14717_ _00571_ net3 mod.u_cpu.rf_ram.memory\[32\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_221_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11929_ _05426_ mod.u_cpu.rf_ram.memory\[221\]\[1\] _05434_ _05436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_127_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11452__I _05106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14648_ _00502_ net3 mod.u_cpu.rf_ram.memory\[363\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_60_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15178__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10068__I _04090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_193_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14579_ _00433_ net3 mod.u_cpu.rf_ram.memory\[398\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_242_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07120_ mod.u_cpu.cpu.bne_or_bge _01429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_70_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__10454__I0 _04423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_158_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08024__A1 _02329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10906__A1 _04732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11954__I0 _05442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10382__A2 _04379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_229_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07953_ mod.u_cpu.rf_ram.memory\[247\]\[0\] _02261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_68_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_229_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_233_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07884_ mod.u_cpu.rf_ram.memory\[221\]\[0\] _02192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_210_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11182__I1 _04658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_255_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_244_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09623_ _03802_ mod.u_cpu.rf_ram.memory\[566\]\[0\] _03830_ _03831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_56_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09554_ _03775_ _03772_ _03776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_83_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07840__I _01482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_224_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08505_ mod.u_cpu.rf_ram.memory\[327\]\[1\] _02812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_58_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09485_ _03704_ _03710_ _03711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_197_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10693__I0 _04579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08436_ mod.u_cpu.rf_ram.memory\[384\]\[1\] mod.u_cpu.rf_ram.memory\[385\]\[1\] mod.u_cpu.rf_ram.memory\[386\]\[1\]
+ mod.u_cpu.rf_ram.memory\[387\]\[1\] _01994_ _02010_ _02743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_168_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_200_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08367_ _02672_ _02673_ _02674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_260_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11398__A1 _04196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_221_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09767__I _03944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_177_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10445__I0 _04410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07318_ _01578_ _01625_ _01626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__14545__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08263__A1 _02523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08298_ _02487_ _02601_ _02604_ _02196_ _02605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_109_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07249_ mod.u_cpu.rf_ram.memory\[477\]\[0\] _01557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__10706__I _04522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12198__I0 mod.u_cpu.rf_ram.memory\[201\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_152_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_178_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10260_ _04250_ _04294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_127_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14695__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_219_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10191_ _04245_ mod.u_cpu.rf_ram.memory\[490\]\[1\] _04243_ _04246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_87_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14114__S _07039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11570__A1 _05187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08620__B _02051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_132_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09208__S _03474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_238_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08318__A2 _02624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13950_ mod.u_arbiter.i_wb_cpu_rdt\[1\] _06906_ _06911_ _03433_ _06924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_74_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12370__I0 _05731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_207_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12901_ _06090_ _01114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_13881_ _06426_ _06670_ _06873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_100_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_234_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2010 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15620_ _01391_ net3 mod.u_cpu.cpu.state.init_done vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_185_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12832_ _06044_ _01091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09451__B _03677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13075__A1 _03713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2021 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_261_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07750__I _01603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2032 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_250_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_215_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2043 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2054 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_215_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15551_ _01322_ net3 mod.u_cpu.cpu.decode.opcode\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2065 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12368__I _03849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_203_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__15320__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12763_ _05998_ mod.u_cpu.rf_ram.memory\[135\]\[1\] _05996_ _05999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_226_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_215_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2076 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2087 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09878__S _04027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14502_ _00356_ net3 mod.u_cpu.rf_ram.memory\[436\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_70_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2098 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_230_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11714_ _05268_ mod.u_cpu.rf_ram.memory\[248\]\[0\] _05285_ _05286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15482_ _01253_ net3 mod.u_arbiter.i_wb_cpu_dbus_adr\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12694_ _05954_ _01043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_203_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14433_ _00287_ net3 mod.u_cpu.rf_ram.memory\[471\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11645_ _05234_ mod.u_cpu.rf_ram.memory\[25\]\[1\] _05236_ _05238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_156_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09677__I _03872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15470__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07688__S0 _01994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14364_ _00218_ net3 mod.u_cpu.rf_ram.memory\[505\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11576_ _04775_ _05191_ _05192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_122_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_171_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13315_ _06412_ _06413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08514__C _01501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10527_ _04467_ mod.u_cpu.rf_ram.memory\[438\]\[1\] _04476_ _04478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_183_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14295_ _00149_ net3 mod.u_cpu.rf_ram.memory\[540\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_109_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12189__I0 _05609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_202_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07197__I _01504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_196_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08006__A1 _02298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_182_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10458_ _04430_ mod.u_cpu.rf_ram.memory\[44\]\[1\] _04427_ _04431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_13246_ _03781_ _06344_ _06348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_237_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11936__I0 mod.u_cpu.rf_ram.memory\[169\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13927__I _06017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09754__A1 _03902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13177_ mod.u_arbiter.i_wb_cpu_rdt\[11\] mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat\[11\]
+ _05781_ _06284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_10389_ _04233_ _04373_ _04385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_83_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12128_ _05422_ _05568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_257_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09506__A1 _01462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12059_ _05521_ mod.u_cpu.rf_ram.memory\[62\]\[0\] _05522_ _05523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_42_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_266_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_237_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_211_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_211_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14418__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_253_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12113__I0 _05550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_244_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_234_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11616__A2 _05130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_206_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_206_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14568__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09270_ _03516_ mod.u_scanchain_local.module_data_in\[43\] _03518_ mod.u_arbiter.i_wb_cpu_dbus_adr\[6\]
+ _03527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_61_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_209_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14015__B1 _06971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08221_ mod.u_cpu.rf_ram.memory\[517\]\[0\] _02529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_53_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_194_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13611__B _03305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12416__I1 _05622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11910__I _05421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13103__S _06234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08152_ _02456_ mod.u_cpu.rf_ram.memory\[548\]\[0\] _02459_ _02460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_158_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08245__A1 _02551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08096__I1 mod.u_cpu.rf_ram.memory\[17\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_158_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10978__I1 _04661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08424__C _02730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_162_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08083_ _01679_ _02391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_88_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_249_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_216_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07835__I _01533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_130_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08985_ mod.u_cpu.cpu.state.o_cnt_r\[1\] mod.u_cpu.cpu.state.o_cnt_r\[0\] mod.u_cpu.cpu.state.o_cnt_r\[3\]
+ mod.u_cpu.cpu.state.o_cnt_r\[2\] _03290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_130_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4907 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4918 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07936_ _01806_ _02244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_151_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4929 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11304__A1 _04868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_229_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_216_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07867_ _02134_ _02175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__15343__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09606_ _03800_ mod.u_cpu.rf_ram.memory\[568\]\[1\] _03815_ _03817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08720__A2 _03023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_56_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_243_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_232_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07798_ _01672_ _02106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__12188__I _05549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09537_ _03760_ _00080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07503__C _01785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_58_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_227_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_212_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_149_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08484__A1 _02041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09468_ _03683_ _03691_ _03694_ _00004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__15493__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_212_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_145_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12280__A2 _05668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_145_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_196_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08419_ _02534_ mod.u_cpu.rf_ram.memory\[412\]\[1\] _02725_ _02726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_212_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09399_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[27\] _03635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09497__I _03722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08615__B _01632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_178_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11430_ _05092_ _00641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_149_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10969__I1 mod.u_cpu.rf_ram.memory\[366\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08334__C _01615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11361_ _03864_ _05047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08787__A2 _03093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13780__A2 _06324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_192_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_256_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11791__A1 _05078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13100_ _06235_ _01168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_10312_ _04168_ _04327_ _04332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_125_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11292_ _05000_ _00595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_14080_ _06904_ mod.u_cpu.rf_ram.memory\[299\]\[1\] _07018_ _07020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_164_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09736__A1 _03902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10243_ _04276_ mod.u_cpu.rf_ram.memory\[482\]\[0\] _04282_ _04283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_13031_ _06186_ mod.u_cpu.rf_ram.memory\[108\]\[0\] _06190_ _06191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_234_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_156_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_156_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12591__I0 _05874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07745__I _01444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_191_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10174_ _04136_ _04234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_117_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_239_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_154_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_266_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_266_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_78_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14982_ _00836_ net3 mod.u_cpu.rf_ram.memory\[213\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_78_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_219_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12343__I0 _05713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_235_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_208_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13933_ _06153_ mod.u_cpu.cpu.bufreg.lsb\[1\] _03390_ _06908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_208_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13048__A1 _06032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13864_ _06856_ _06857_ _01310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_19_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14710__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07480__I _01787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14096__I0 _07021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_235_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15603_ _01374_ net3 mod.u_cpu.rf_ram.memory\[117\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08509__C _02677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12815_ _02317_ _06031_ _06033_ _01085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_16_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07413__C _01720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13795_ _06331_ _06794_ _06795_ _06735_ _06796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_90_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_203_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09511__I1 _03735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15534_ _01305_ net3 mod.u_cpu.cpu.immdec.imm30_25\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_43_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12746_ _05984_ mod.u_cpu.rf_ram.memory\[219\]\[1\] _05986_ _05988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08475__A1 _02022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_203_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10282__A1 _04311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14860__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_175_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15465_ _01239_ net3 mod.u_cpu.cpu.ctrl.o_ibus_adr\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12677_ _05938_ mod.u_cpu.rf_ram.memory\[143\]\[1\] _05941_ _05943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_129_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14416_ _00270_ net3 mod.u_cpu.rf_ram.memory\[47\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11628_ _04106_ _05226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__13220__A1 _06122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15396_ _01171_ net3 mod.u_cpu.rf_ram.memory\[101\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_128_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_156_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09975__A1 _03714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_200_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13771__A2 _06772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14347_ _00201_ net3 mod.u_cpu.rf_ram.memory\[514\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11559_ _05047_ _05171_ _05181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_183_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15216__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14278_ _00132_ net3 mod.u_cpu.rf_ram.memory\[548\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_171_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13229_ mod.u_arbiter.i_wb_cpu_rdt\[30\] _03456_ _06335_ _06336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_143_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08086__S0 _02349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_170_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07655__I _01644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_97_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_170_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14240__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15366__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08770_ _02293_ _03069_ _03076_ _02321_ _03077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12334__I0 _05696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07721_ _02027_ _02028_ _02029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08702__A2 _03000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12002__S _05481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07652_ _01749_ _01960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_38_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14390__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_225_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_214_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_214_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_207_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07583_ _01890_ _01891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_20_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12637__I1 mod.u_cpu.rf_ram.memory\[148\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_209_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09322_ _03542_ _03538_ _03570_ _03559_ _03571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XANTENNA__08466__A1 _01864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_222_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_221_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09253_ _03479_ mod.u_scanchain_local.module_data_in\[40\] _03408_ mod.u_arbiter.i_wb_cpu_dbus_adr\[3\]
+ _03513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_181_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_222_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08204_ _02478_ mod.u_cpu.rf_ram.memory\[564\]\[0\] _02511_ _02512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_194_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09184_ _03463_ _00021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_182_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13062__I1 _06005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08135_ _02150_ _02435_ _02442_ _02185_ _02443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_175_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08313__S1 _02454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13762__A2 mod.u_cpu.cpu.immdec.imm24_20\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_257_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08066_ _01823_ _02373_ _02374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_31_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10820__I0 _04666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_257_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09718__A1 _03902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_255_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10328__A2 _03886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11087__I _03780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_248_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13278__A1 _06306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08968_ mod.u_arbiter.i_wb_cpu_dbus_we _03263_ mod.u_cpu.cpu.immdec.imm24_20\[0\]
+ _03273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_102_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14733__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13278__B2 _06372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12325__I0 _05692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07919_ _02070_ mod.u_cpu.rf_ram.memory\[212\]\[0\] _02227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_57_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11828__A2 _05362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08899_ _02039_ _03186_ _03205_ _03206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_84_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11815__I _03949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10930_ _04749_ _04733_ _04750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__14078__I0 _06578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_264_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07752__I0 mod.u_cpu.rf_ram.memory\[148\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14883__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10861_ _04702_ _04703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_260_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12600_ _05891_ mod.u_cpu.rf_ram.memory\[155\]\[1\] _05889_ _05892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XPHY_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_213_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13580_ _06610_ _01273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10792_ _04637_ mod.u_cpu.rf_ram.memory\[394\]\[0\] _04655_ _04656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_213_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08847__I3 mod.u_cpu.rf_ram.memory\[35\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_12531_ _05593_ _04528_ _05846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XPHY_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_235_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_184_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_200_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08345__B _02651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__15239__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_15250_ _00075_ net4 mod.u_arbiter.i_wb_cpu_rdt\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_185_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12462_ mod.u_arbiter.i_wb_cpu_ack _03406_ _05800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_240_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_200_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_200_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_200_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14201_ _06152_ _06151_ _06056_ _07097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_11413_ _05081_ _00635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09957__A1 _03905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13753__A2 _06472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15181_ _01034_ net3 mod.u_cpu.rf_ram.memory\[144\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12393_ _01609_ _05747_ _05748_ _00948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__11764__A1 _04227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_197_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14132_ _03850_ _05631_ _07053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_32_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11344_ _05035_ _00612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__14263__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15389__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14063_ mod.u_arbiter.i_wb_cpu_rdt\[29\] _06937_ _07004_ mod.u_arbiter.i_wb_cpu_dbus_dat\[29\]
+ _07009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_4_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11275_ _04987_ _00591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_165_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10319__A2 _04336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12564__I0 _05855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09024__I3 mod.u_arbiter.i_wb_cpu_dbus_dat\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13014_ _06179_ _01138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_10226_ mod.u_cpu.rf_ram.memory\[485\]\[1\] _04111_ _04269_ _04271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_10157_ _04220_ _00240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_66_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14965_ _00819_ net3 mod.u_cpu.rf_ram.memory\[569\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10088_ _04157_ mod.u_cpu.rf_ram.memory\[504\]\[1\] _04169_ _04171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_208_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11725__I _03857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13916_ _06894_ _06895_ _01324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_48_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08696__A1 _03001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14896_ _00750_ net3 mod.u_cpu.rf_ram.memory\[236\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_207_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_262_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_165_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13847_ _06803_ _06841_ _06842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_90_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13816__I0 mod.u_arbiter.i_wb_cpu_rdt\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12757__S _05993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_250_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13778_ _06404_ _06744_ _06779_ _06426_ _06780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_203_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10255__A1 _04290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15517_ _01288_ net3 mod.u_cpu.rf_ram.memory\[309\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_149_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12729_ _05966_ mod.u_cpu.rf_ram.memory\[78\]\[1\] _05975_ _05977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_241_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_175_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15448_ _01222_ net3 mod.u_cpu.cpu.ctrl.o_ibus_adr\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_175_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14606__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13744__A2 _06139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_191_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15379_ _01154_ net3 mod.u_cpu.rf_ram.memory\[69\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_156_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_209_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08620__A1 _02046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_239_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_172_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08702__C _02852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12291__I _05604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09940_ _04044_ _04069_ _04070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_125_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14756__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09871_ _04018_ mod.u_cpu.rf_ram.memory\[538\]\[1\] _04020_ _04022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_217_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_258_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08822_ _02405_ _03125_ _03128_ _02415_ _03129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10030__I1 mod.u_cpu.rf_ram.memory\[512\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10730__A2 _04599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13336__B _06432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08753_ mod.u_cpu.rf_ram.memory\[101\]\[1\] _03060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_61_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_254_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07704_ mod.u_cpu.rf_ram.memory\[261\]\[0\] _02012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_54_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14011__I _06970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08684_ _02230_ _02990_ _02991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_66_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_227_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13680__A1 _06689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09105__I net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07635_ _01915_ _01933_ _01942_ _01768_ _01943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_1908 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08782__S1 _02107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_253_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13807__I0 mod.u_arbiter.i_wb_cpu_rdt\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_242_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12235__A2 _05640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07566_ _01665_ _01874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_263_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14167__B _07076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_181_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09305_ _03554_ mod.u_scanchain_local.module_data_in\[49\] _03555_ mod.u_arbiter.i_wb_cpu_dbus_adr\[12\]
+ _03556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_94_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_210_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11294__I0 _04978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_224_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_194_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13983__A2 _06938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07497_ _01517_ mod.u_cpu.rf_ram.memory\[444\]\[0\] _01804_ _01805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10797__A2 _04644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09976__S _04093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09236_ _03414_ _03400_ _03497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_194_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14286__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09939__A1 _04033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13735__A2 _03424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_181_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15531__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09167_ _03453_ _00013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_175_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11746__A1 _02412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12794__I0 _06019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09775__I _03950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08118_ mod.u_cpu.rf_ram.memory\[32\]\[0\] mod.u_cpu.rf_ram.memory\[33\]\[0\] mod.u_cpu.rf_ram.memory\[34\]\[0\]
+ mod.u_cpu.rf_ram.memory\[35\]\[0\] _02403_ _02383_ _02426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_266_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_181_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__08611__A1 _02074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09098_ _03398_ mod.u_cpu.cpu.state.ibus_cyc _03399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_163_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_79_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08049_ mod.u_cpu.rf_ram.memory\[71\]\[0\] _02357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_162_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11060_ _04827_ mod.u_cpu.rf_ram.memory\[352\]\[0\] _04839_ _04840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_135_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_192_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10011_ _04050_ _04117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_5224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_114_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_249_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_130_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_105 la_data_out[23] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_5257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xtiny_user_project_116 la_data_out[34] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_127 la_data_out[45] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_5268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_138 la_data_out[56] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_3800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_185_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xtiny_user_project_149 wbs_ack_o vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__11545__I _05124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_218_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14750_ _00604_ net3 mod.u_cpu.rf_ram.memory\[312\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08678__A1 _02543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11962_ _05458_ _00807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12474__A2 _04033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_244_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09015__I mod.u_cpu.cpu.state.o_cnt_r\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13701_ mod.u_cpu.cpu.immdec.imm19_12_20\[3\] _06708_ _06709_ _06710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_3877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_151_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10913_ _01880_ _04737_ _04738_ _00478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_3888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14681_ _00535_ net3 mod.u_cpu.rf_ram.memory\[347\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11893_ _05410_ _00786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3899 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_232_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15061__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13632_ _06319_ _06324_ _06643_ _06644_ _06645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_71_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10844_ _04690_ _00457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07898__C _02049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_164_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_201_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14629__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13563_ mod.u_arbiter.i_wb_cpu_dbus_adr\[15\] mod.u_arbiter.i_wb_cpu_dbus_adr\[16\]
+ _06599_ _06601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_185_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10775_ _04643_ _04644_ _04645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_201_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15302_ _00062_ net4 mod.u_scanchain_local.module_data_in\[59\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_157_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12514_ _05395_ _05667_ _05835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_160_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08850__A1 _02356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13494_ _03631_ _06551_ _06552_ _03635_ _06555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_173_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_205_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_201_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15233_ _01086_ net3 mod.u_cpu.rf_ram.memory\[127\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_185_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12445_ _05782_ _05783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_139_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__14779__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09685__I _03822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08602__A1 _01852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15164_ _01017_ net3 mod.u_cpu.rf_ram.memory\[152\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_176_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12376_ _05737_ _00942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_165_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_197_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14115_ _07042_ _01376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_11327_ _05014_ mod.u_cpu.rf_ram.memory\[311\]\[1\] _05021_ _05024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_181_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15095_ _00949_ net3 mod.u_cpu.rf_ram.memory\[509\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_125_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_153_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10960__A2 _04713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14046_ _06995_ _06996_ _01353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_141_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11258_ _04975_ _00586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_141_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13935__I _06909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_1243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_136_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10209_ _03942_ _04173_ _04259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_95_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11189_ _04928_ _00564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_67_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08461__S0 _01837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14948_ _00802_ net3 mod.u_cpu.rf_ram.memory\[21\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08669__A1 _02711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15404__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13662__A1 _06434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_236_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_263_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_224_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10476__A1 _04299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_235_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14879_ _00733_ net3 mod.u_cpu.rf_ram.memory\[248\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_1_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_224_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07341__A1 _01647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07420_ _01604_ _01728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_165_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_251_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07892__A2 mod.u_cpu.rf_ram.memory\[218\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_189_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_245_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_206_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08516__S1 _02748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07351_ mod.u_cpu.raddr\[2\] _01659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__15554__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07282_ _01486_ _01554_ _01589_ _01590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_137_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_206_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09021_ _03298_ _03255_ _03326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_191_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13717__A2 mod.u_arbiter.i_wb_cpu_rdt\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09641__I0 _03802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08432__C _01918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09923_ _04054_ mod.u_cpu.rf_ram.memory\[530\]\[1\] _04056_ _04058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_252_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12153__A1 _05312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_259_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_213_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10003__I1 _04111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09854_ _03782_ _04003_ _04010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_24_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08805_ _02063_ _03108_ _03111_ _01669_ _03112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09785_ _03957_ _00131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_46_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11365__I _05031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07580__A1 _01872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08736_ mod.u_cpu.rf_ram.memory\[255\]\[1\] _03043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_73_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15084__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13653__A1 _06447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_226_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__12700__I0 _05938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_227_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_199_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08667_ mod.u_cpu.rf_ram.memory\[217\]\[1\] _02974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_1705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_214_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07618_ mod.u_cpu.rf_ram.memory\[319\]\[0\] _01926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08598_ mod.u_cpu.rf_ram.memory\[263\]\[1\] _02905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_183_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_241_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_198_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07549_ _01856_ _01857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_224_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07635__A2 _01933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08832__A1 _02150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10560_ _04209_ _04487_ _04500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__14921__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_220_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09880__I0 _04018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_210_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09219_ mod.u_arbiter.i_wb_cpu_dbus_dat\[31\] _03483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_194_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10491_ _04453_ mod.u_cpu.rf_ram.memory\[444\]\[0\] _04454_ _04455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_120_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_12230_ _05322_ _05637_ _05638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_136_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07399__A1 _01567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12392__A1 _05581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12161_ mod.u_cpu.rf_ram.memory\[73\]\[0\] _05437_ _05590_ _05591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_163_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08691__S0 _02349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_190_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11112_ _04876_ _00539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_1_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12092_ _05408_ _05543_ _05544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_150_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_235_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xtiny_user_project_11 io_oeb[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_77_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5010 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11043_ _04827_ mod.u_cpu.rf_ram.memory\[355\]\[0\] _04828_ _04829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_104_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5021 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08899__A1 _02039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtiny_user_project_22 io_oeb[14] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_5032 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14301__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13892__A1 _03872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_33 io_oeb[25] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__15427__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtiny_user_project_44 io_oeb[36] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_5043 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_118_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xtiny_user_project_55 io_out[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_5054 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xtiny_user_project_66 io_out[22] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_5065 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5076 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_77 io_out[33] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_92_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5087 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_77_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_88 la_data_out[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_99 la_data_out[17] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_5098 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14802_ _00656_ net3 mod.u_cpu.rf_ram.memory\[286\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_4353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12994_ _06165_ _01132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_4386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_264_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_245_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14733_ _00587_ net3 mod.u_cpu.rf_ram.memory\[321\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11945_ _04983_ _03837_ _05447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_166_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14451__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_217_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_206_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15577__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2940 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2951 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2962 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_233_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14664_ _00518_ net3 mod.u_cpu.rf_ram.memory\[355\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2973 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07874__A2 _02181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11876_ _05395_ _05397_ _05398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2984 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2995 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13615_ _04844_ _05020_ _06633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10619__I _03773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10827_ _04621_ _04679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_14595_ _00449_ net3 mod.u_cpu.rf_ram.memory\[390\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_242_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11958__A1 _05047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_203_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13546_ _06591_ _01258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08823__A1 _02365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10758_ _04626_ mod.u_cpu.rf_ram.memory\[400\]\[1\] _04631_ _04633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09871__I0 _04018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10630__A1 _04412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_200_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13477_ _06544_ _01236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_145_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10689_ _04587_ _00405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_15216_ _01069_ net3 mod.u_cpu.rf_ram.memory\[134\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_103_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_145_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12428_ _05759_ _05771_ _05772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__09623__I0 _03802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10354__I _03865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15147_ _01000_ net3 mod.u_cpu.rf_ram.memory\[161\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_153_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12359_ _05666_ _05725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_153_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_15078_ _00932_ net3 mod.u_cpu.rf_ram.memory\[182\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_114_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_206_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_253_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14029_ mod.u_arbiter.i_wb_cpu_dbus_dat\[21\] _06978_ _06984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09926__I1 mod.u_cpu.rf_ram.memory\[52\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12686__A2 _05947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13883__A1 _06468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09570_ _03787_ _03788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_23_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_83_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_208_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08521_ _01893_ mod.u_cpu.rf_ram.memory\[340\]\[1\] _02827_ _02828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_236_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_224_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_224_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08452_ _01615_ _02759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_91_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14944__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_212_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07403_ _01710_ _01711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_223_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_196_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13938__A2 _06909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08383_ _02687_ _02689_ _02077_ _02690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09067__A1 _03353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14060__A1 mod.u_arbiter.i_wb_cpu_rdt\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08114__I0 mod.u_cpu.rf_ram.memory\[48\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_149_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_220_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07334_ _01607_ mod.u_cpu.rf_ram.memory\[492\]\[0\] _01641_ _01642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09862__I0 _04001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10621__A1 _04542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07265_ _01510_ _01573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_149_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09004_ _03303_ _03309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07196_ _01503_ _01504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_219_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_192_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12374__A1 _05563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08162__C _02469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_145_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14324__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09790__A2 _03961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13174__I0 mod.u_arbiter.i_wb_cpu_rdt\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09906_ _04046_ _00163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_59_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_263_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_150_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13874__A1 _06412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12921__I0 _06088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_258_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09837_ _02576_ _03997_ _03998_ _00142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_59_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14474__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07553__A1 _01857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_230_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09768_ _03945_ _03943_ _03946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_246_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_227_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08719_ _02751_ mod.u_cpu.rf_ram.memory\[230\]\[1\] _03025_ _02154_ _03026_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_227_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09699_ _03889_ _03890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_132_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07305__A1 _01578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_70_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11730_ _05296_ _00737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_215_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_2269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_265_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_202_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13229__I1 _03456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11661_ _05248_ _00716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_186_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07241__C _01529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09058__A1 _03306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_199_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_186_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13400_ _06434_ _06494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_168_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10612_ _04523_ mod.u_cpu.rf_ram.memory\[424\]\[0\] _04535_ _04536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08805__A1 _02063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14380_ _00234_ net3 mod.u_cpu.rf_ram.memory\[497\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11592_ _05202_ _00693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_167_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13331_ _06424_ _06370_ _06427_ _06417_ _06428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_70_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11660__I0 _05243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10543_ _04486_ mod.u_cpu.rf_ram.memory\[435\]\[0\] _04488_ _04489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08900__S1 _02495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08281__A2 mod.u_cpu.rf_ram.memory\[460\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09449__B _03677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13262_ _05782_ mod.u_arbiter.i_wb_cpu_rdt\[7\] _06360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_143_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10474_ _04435_ _04442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_15001_ _00855_ net3 mod.u_cpu.rf_ram.memory\[67\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11168__A2 _04906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12213_ _05625_ _00891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_108_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10174__I _04136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13193_ _06299_ _06300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_159_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12144_ _05566_ mod.u_cpu.rf_ram.memory\[75\]\[1\] _05577_ _05579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_151_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09781__A2 _03829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14817__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07792__A1 _02097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13165__I0 _06273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09908__I1 mod.u_cpu.rf_ram.memory\[532\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12075_ _05532_ _00846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_173_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08416__S0 _02225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13865__A1 _06282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11026_ _04412_ _04780_ _04816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_133_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10679__A1 _04307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11934__S _05439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14967__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11479__I0 _05114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09297__A1 mod.u_cpu.cpu.ctrl.o_ibus_adr\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12977_ _03269_ _06152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13093__A2 _03878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_206_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13632__A4 _06644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11928_ _02192_ _05434_ _05435_ _00796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_14716_ _00570_ net3 mod.u_cpu.rf_ram.memory\[32\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10151__I0 _04215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_233_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09203__I _03414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_205_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14647_ _00501_ net3 mod.u_cpu.rf_ram.memory\[364\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_260_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11859_ _05310_ _05385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_162_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14042__A1 mod.u_arbiter.i_wb_cpu_rdt\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_221_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_202_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_202_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_193_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13396__A3 _06490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14578_ _00432_ net3 mod.u_cpu.rf_ram.memory\[398\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_192_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_186_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10603__A1 _04527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11651__I0 _05234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10454__I1 mod.u_cpu.rf_ram.memory\[44\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13529_ _06236_ _06581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_118_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_203_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10285__S _04310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14347__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_146_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_174_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10084__I _03804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09873__I _03915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11954__I1 mod.u_cpu.rf_ram.memory\[218\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_217_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14497__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07952_ _02175_ mod.u_cpu.rf_ram.memory\[244\]\[0\] _02259_ _02260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_141_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13856__A1 _06397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07393__I _01700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_233_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_68_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_229_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07883_ _02190_ _02191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_29_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09622_ _03814_ _03829_ _03830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_95_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_256_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_249_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14220__S _07106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10390__I0 _04365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_228_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_209_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_209_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09553_ _03774_ _03775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_83_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08504_ _02041_ mod.u_cpu.rf_ram.memory\[324\]\[1\] _02810_ _02811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11095__A1 _04457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_224_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09484_ _03707_ _03709_ _03710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__07838__A2 _02145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_252_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_211_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08435_ _02609_ _02732_ _02741_ _02742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__15122__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_197_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__12675__S _05941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08366_ mod.u_cpu.rf_ram.memory\[487\]\[1\] _02673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__08952__I _03256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08638__I1 mod.u_cpu.rf_ram.memory\[169\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_177_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11398__A2 _03975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13792__B1 _06402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10445__I1 mod.u_cpu.rf_ram.memory\[451\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07317_ mod.u_cpu.rf_ram.memory\[487\]\[0\] _01625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_192_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08263__A2 _02562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08297_ _02191_ mod.u_cpu.rf_ram.memory\[454\]\[1\] _02603_ _02093_ _02604_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_109_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15272__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07248_ _01539_ _01556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_191_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12347__A1 _04014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12198__I1 _05437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07179_ _01419_ _01443_ _01487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_11_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_191_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10190_ _04177_ _04245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_156_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07774__A1 _02080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11570__A2 _05130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_259_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_235_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12370__I1 mod.u_cpu.rf_ram.memory\[499\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12900_ _06088_ mod.u_cpu.rf_ram.memory\[96\]\[0\] _06089_ _06090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_19_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_262_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13880_ _06811_ _06871_ _06872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_143_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_235_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12831_ _06035_ mod.u_cpu.rf_ram.memory\[124\]\[0\] _06043_ _06044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_2000 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_189_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_62_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2011 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09279__A1 mod.u_cpu.cpu.ctrl.o_ibus_adr\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_265_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13075__A2 _05640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2022 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2033 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15550_ _01321_ net3 mod.u_cpu.cpu.csr_d_sel vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_43_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2044 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_203_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2055 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12762_ _05937_ _05998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2066 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2077 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14501_ _00355_ net3 mod.u_cpu.rf_ram.memory\[437\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2088 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11713_ _05283_ _05284_ _05285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_203_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08067__C _02359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15481_ _00004_ net3 mod.u_cpu.cpu.bufreg.c_r vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2099 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_242_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_187_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12693_ mod.u_cpu.rf_ram.memory\[141\]\[0\] _05622_ _05953_ _05954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14432_ _00286_ net3 mod.u_cpu.rf_ram.memory\[471\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11644_ _05237_ _00710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_204_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15615__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14363_ _00217_ net3 mod.u_cpu.rf_ram.memory\[506\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11575_ _05119_ _05191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07688__S1 _01995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_196_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_183_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13314_ _06138_ _06412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_6_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10526_ _04477_ _00352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_182_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14294_ _00148_ net3 mod.u_cpu.rf_ram.memory\[540\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_13_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_171_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11929__S _05434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13245_ _06347_ _01201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_109_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10457_ _04429_ _04430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_108_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09693__I _03884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11936__I1 _05230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09754__A2 _03933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13176_ _06282_ _06283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_124_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10388_ _04384_ _00307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_170_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12127_ _05567_ _00863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_151_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13838__A1 _03331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09506__A2 mod.u_cpu.rf_ram_if.wdata1_r\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08102__I _01646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12058_ _05428_ _03878_ _05522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_77_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_250_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07146__C _01425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11009_ _04804_ _04788_ _04805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_238_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07941__I _01539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_252_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08190__A1 _02457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15145__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_206_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12113__I1 mod.u_cpu.rf_ram.memory\[68\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11077__A1 _04852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_240_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10124__I0 _04193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_221_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07376__S0 _01682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14015__A1 mod.u_arbiter.i_wb_cpu_rdt\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14015__B2 mod.u_arbiter.i_wb_cpu_dbus_dat\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_221_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_221_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15295__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08220_ _01538_ _02528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_166_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_221_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12577__A1 _05428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11624__I0 _05222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_193_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08151_ _02457_ _02458_ _02459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_159_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09442__A1 _03663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08245__A2 _02552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10807__I _04640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_186_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07388__I _01695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_174_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_146_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08082_ mod.u_cpu.rf_ram.memory\[8\]\[0\] mod.u_cpu.rf_ram.memory\[9\]\[0\] mod.u_cpu.rf_ram.memory\[10\]\[0\]
+ mod.u_cpu.rf_ram.memory\[11\]\[0\] _02171_ _02267_ _02390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_179_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11001__A1 _04527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_142_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08984_ _03286_ _03287_ _03288_ _01421_ _03289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XANTENNA__09108__I _03407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4908 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07935_ mod.u_cpu.rf_ram.memory\[232\]\[0\] mod.u_cpu.rf_ram.memory\[233\]\[0\] mod.u_cpu.rf_ram.memory\[234\]\[0\]
+ mod.u_cpu.rf_ram.memory\[235\]\[0\] _02242_ _02172_ _02243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_4919 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_244_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07866_ _02154_ _02174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_56_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08947__I _03251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_257_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10363__I0 _04365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_35 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09605_ _03816_ _00092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_186_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_28_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07797_ _01488_ _02105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09536_ _03740_ mod.u_cpu.rf_ram.memory\[574\]\[0\] _03759_ _03760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_58_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10115__I0 _04162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14512__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15638__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_197_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_197_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_184_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_224_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_184_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09467_ _03693_ _03694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08484__A2 mod.u_cpu.rf_ram.memory\[356\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_223_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_185_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08418_ _02526_ _02724_ _02725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_145_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_212_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_200_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09398_ _03632_ _03633_ _03634_ _00068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_184_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14662__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08349_ _01841_ _02656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_165_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11360_ _05045_ _05046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_164_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11791__A2 _05320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10311_ _04331_ _00283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_11291_ _04999_ mod.u_cpu.rf_ram.memory\[317\]\[1\] _04997_ _05000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08619__S0 _02066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15018__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13030_ _03904_ _06092_ _06190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12040__I0 _05498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09736__A2 _03919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10242_ _04281_ _04263_ _04282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_3_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_191_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_65_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10173_ _03904_ _04233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_121_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15168__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14981_ _00835_ net3 mod.u_cpu.rf_ram.memory\[60\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_43_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13932_ _03268_ mod.u_cpu.cpu.bufreg.lsb\[1\] _03279_ _03269_ _06907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_120_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_263_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_232_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_234_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13863_ mod.u_cpu.cpu.immdec.imm24_20\[2\] _06836_ _06837_ mod.u_cpu.cpu.immdec.imm24_20\[3\]
+ _06857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__13048__A2 _06201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_250_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11059__A1 _04838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15602_ _01373_ net3 mod.u_cpu.rf_ram.memory\[117\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12814_ _06032_ _06031_ _06033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_222_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13794_ _06726_ _06407_ _06486_ _06795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_188_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11854__I0 _05366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12745_ _02199_ _05986_ _05987_ _01061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_15533_ _01304_ net3 mod.u_cpu.cpu.immdec.imm30_25\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10282__A2 _04310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15464_ _01238_ net3 mod.u_cpu.cpu.ctrl.o_ibus_adr\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12676_ _05942_ _01037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_203_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14415_ _00269_ net3 mod.u_cpu.rf_ram.memory\[480\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_8_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11627_ _05225_ _00705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_15395_ _01170_ net3 mod.u_cpu.rf_ram.memory\[101\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_128_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13220__A2 _06123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10034__A2 _03665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_14346_ _00200_ net3 mod.u_cpu.rf_ram.memory\[514\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11558_ _05143_ _05180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_200_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09975__A2 _04077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10509_ _04466_ _00346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_14277_ _00131_ net3 mod.u_cpu.rf_ram.memory\[54\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11489_ _01999_ _05131_ _05134_ _00658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_170_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13228_ _06334_ _06335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_174_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08086__S1 _02393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08786__I0 mod.u_cpu.rf_ram.memory\[88\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13159_ mod.u_arbiter.i_wb_cpu_rdt\[30\] mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat\[14\]
+ _06268_ _06271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_257_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_214_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_250_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07720_ mod.u_cpu.rf_ram.memory\[271\]\[0\] _02028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_211_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11298__A1 _04457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_239_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10345__I0 _04348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14535__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07671__I _01914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_253_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07651_ mod.u_cpu.rf_ram.memory\[296\]\[0\] mod.u_cpu.rf_ram.memory\[297\]\[0\] mod.u_cpu.rf_ram.memory\[298\]\[0\]
+ mod.u_cpu.rf_ram.memory\[299\]\[0\] _01957_ _01958_ _01959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_168_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12098__I0 _05539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07582_ _01487_ _01890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_53_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_207_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_241_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_209_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09321_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[11\] mod.u_cpu.cpu.ctrl.o_ibus_adr\[10\] _03570_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_179_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14685__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_222_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_206_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_209_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09252_ _03507_ _03511_ _03512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_209_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_167_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_261_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08203_ _02509_ _02510_ _02511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09183_ mod.u_arbiter.i_wb_cpu_rdt\[18\] mod.u_arbiter.i_wb_cpu_dbus_dat\[15\] _03459_
+ _03463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_08134_ _02155_ _02438_ _02441_ _02166_ _02442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__12270__I0 _05660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_179_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07521__S0 _01826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_179_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08065_ mod.u_cpu.rf_ram.memory\[79\]\[0\] _02373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_146_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07846__I _01749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_190_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09718__A2 _03905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_216_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07729__A1 _01471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15310__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_249_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_192_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_130_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08967_ mod.u_arbiter.i_wb_cpu_dbus_we _03271_ _03263_ _03272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XTAP_4705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07918_ mod.u_cpu.rf_ram.memory\[213\]\[0\] _02226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_116_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_245_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08898_ _03195_ _03204_ _02520_ _03205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_57_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_216_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15460__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_217_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07849_ _01681_ _02157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_57_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14078__I1 mod.u_cpu.rf_ram.memory\[299\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_232_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_186_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_232_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12089__I0 _05533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10860_ _03992_ _04134_ _04701_ _04702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_204_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_227_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09519_ _03703_ _03742_ _03743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XPHY_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_231_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12927__I _06072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10791_ _04242_ _04648_ _04655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_197_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_73_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12530_ _05845_ _00988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_213_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_262_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07760__S0 _02066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08345__C _02377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12461_ _03359_ _03355_ _05798_ _05799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__10447__I _04347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_228_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_166_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14200_ _06046_ _06151_ _07096_ _01408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_11412_ mod.u_cpu.rf_ram.memory\[297\]\[1\] _05065_ _05079_ _05081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_15180_ _01033_ net3 mod.u_cpu.rf_ram.memory\[144\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_165_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12392_ _05581_ _05747_ _05748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_201_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_201_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07968__A1 _02174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14408__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_181_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14131_ _07052_ _01382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11764__A2 _05319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11343_ _05028_ mod.u_cpu.rf_ram.memory\[308\]\[0\] _05034_ _05035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_165_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_193_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14062_ mod.u_arbiter.i_wb_cpu_dbus_dat\[30\] _07000_ _07008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_10_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11274_ _04976_ mod.u_cpu.rf_ram.memory\[31\]\[1\] _04985_ _04987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_234_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11278__I _04989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13013_ _06107_ mod.u_cpu.rf_ram.memory\[85\]\[0\] _06178_ _06179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_10225_ _01622_ _04269_ _04270_ _00258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_152_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10575__I0 _04498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14558__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_239_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09971__I _03762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08393__A1 _02083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10156_ _04217_ mod.u_cpu.rf_ram.memory\[494\]\[0\] _04219_ _04220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_67_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_208_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_208_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14964_ _00818_ net3 mod.u_cpu.rf_ram.memory\[569\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10087_ _04170_ _00220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_181_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_235_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13915_ _05790_ _06413_ _06811_ _06465_ _06895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__08535__I3 mod.u_cpu.rf_ram.memory\[299\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14895_ _00749_ net3 mod.u_cpu.rf_ram.memory\[237\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_78_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_251_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_223_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13846_ _06437_ _06662_ _06840_ _06841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_223_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13816__I1 mod.u_arbiter.i_wb_cpu_rdt\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13777_ _06667_ _06778_ _06779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__11741__I _05249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_188_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10989_ _04790_ _00502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_43_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08536__B _02207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15516_ _01287_ net3 mod.u_cpu.rf_ram.memory\[319\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_15_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10255__A2 _04137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_206_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12728_ _05976_ _01055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_31_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12659_ _05930_ _01032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_15447_ _01221_ net3 mod.u_cpu.cpu.ctrl.o_ibus_adr\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_129_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12252__I0 _05635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_15378_ _01153_ net3 mod.u_cpu.rf_ram.memory\[82\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_129_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15333__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14329_ _00183_ net3 mod.u_cpu.rf_ram.memory\[523\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08620__A2 _02926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_143_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_217_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09870_ _04021_ _00152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15483__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_225_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08821_ _02410_ mod.u_cpu.rf_ram.memory\[30\]\[1\] _03127_ _01830_ _03128_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_239_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08752_ mod.u_cpu.rf_ram.memory\[96\]\[1\] mod.u_cpu.rf_ram.memory\[97\]\[1\] mod.u_cpu.rf_ram.memory\[98\]\[1\]
+ mod.u_cpu.rf_ram.memory\[99\]\[1\] _02211_ _02386_ _03059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_227_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08136__A1 _02149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07703_ mod.u_cpu.rf_ram.memory\[256\]\[0\] mod.u_cpu.rf_ram.memory\[257\]\[0\] mod.u_cpu.rf_ram.memory\[258\]\[0\]
+ mod.u_cpu.rf_ram.memory\[259\]\[0\] _01994_ _02010_ _02011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_2_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_227_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08683_ _02594_ _02986_ _02989_ _02591_ _02990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_66_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_93_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_214_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07634_ _01918_ _01937_ _01941_ _01929_ _01942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_1909 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_246_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13807__I1 mod.u_arbiter.i_wb_cpu_rdt\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_213_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07565_ mod.u_cpu.rf_ram.memory\[368\]\[0\] mod.u_cpu.rf_ram.memory\[369\]\[0\] mod.u_cpu.rf_ram.memory\[370\]\[0\]
+ mod.u_cpu.rf_ram.memory\[371\]\[0\] _01843_ _01844_ _01873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__08439__A2 _02745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_224_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_210_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09304_ _03407_ _03555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_179_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_222_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11294__I1 mod.u_cpu.rf_ram.memory\[316\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07496_ _01802_ _01803_ _01804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_179_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_224_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_194_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07742__S0 _02048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_181_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09235_ _03495_ _03496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_194_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10267__I _03751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_210_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_166_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_194_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09166_ mod.u_arbiter.i_wb_cpu_rdt\[11\] mod.u_arbiter.i_wb_cpu_dbus_dat\[8\] _03452_
+ _03453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_33_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09939__A2 _04068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13578__I _03692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11746__A2 _05306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12943__A1 _05784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08117_ _02420_ _02422_ _02423_ _02424_ _02391_ _01552_ _02425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__08998__I0 _03276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_257_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09097_ net5 _03398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_174_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08611__A2 _02917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_266_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14700__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08048_ _01993_ _02356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_150_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_192_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10010_ _04116_ _00197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_5214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_89_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_130_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_130_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09999_ _04077_ _04108_ _04109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_5247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_106 la_data_out[24] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_103_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14850__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13019__S _06182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtiny_user_project_117 la_data_out[35] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_5258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_130_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xtiny_user_project_128 la_data_out[46] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_264_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xtiny_user_project_139 la_data_out[57] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_4535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_217_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13120__A1 _03941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09324__B1 _03402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_4568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11961_ _05450_ mod.u_cpu.rf_ram.memory\[529\]\[1\] _05456_ _05458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_91_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08678__A2 _02981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_178_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_217_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_56_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_233_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13700_ _06655_ _06709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_10912_ _04611_ _04737_ _04738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__11682__A1 _04700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14680_ _00534_ net3 mod.u_cpu.rf_ram.memory\[347\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__15206__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11892_ _05385_ mod.u_cpu.rf_ram.memory\[226\]\[0\] _05409_ _05410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_205_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_260_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13631_ _06371_ _06310_ _06644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_72_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10843_ _04682_ mod.u_cpu.rf_ram.memory\[386\]\[1\] _04688_ _04690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_44_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_220_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_25_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_198_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08356__B _01618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_73_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13562_ _06600_ _01265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_197_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10774_ _03723_ _04225_ _04644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__12482__I0 _05813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_198_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_200_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__14230__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12513_ _05834_ _00982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_13_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15301_ _00061_ net4 mod.u_scanchain_local.module_data_in\[58\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_185_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15356__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_197_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13493_ _06554_ _01242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__08850__A2 mod.u_cpu.rf_ram.memory\[36\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_185_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12444_ _05781_ _05782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_15232_ _01085_ net3 mod.u_cpu.rf_ram.memory\[127\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_138_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13488__I _06537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15163_ _01016_ net3 mod.u_cpu.rf_ram.memory\[153\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12375_ _05731_ mod.u_cpu.rf_ram.memory\[17\]\[0\] _05736_ _05737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_126_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10905__I _04708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08602__A2 _02901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_154_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11002__S _04799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14380__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14114_ _07041_ mod.u_cpu.rf_ram.memory\[87\]\[1\] _07039_ _07042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_114_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11326_ _01939_ _05021_ _05023_ _00606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_125_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15094_ _00948_ net3 mod.u_cpu.rf_ram.memory\[509\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_158_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14045_ mod.u_arbiter.i_wb_cpu_rdt\[24\] _06987_ _06993_ mod.u_arbiter.i_wb_cpu_dbus_dat\[24\]
+ _06996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_141_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11257_ _04961_ mod.u_cpu.rf_ram.memory\[321\]\[0\] _04974_ _04975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_158_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10841__S _04688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10208_ _04258_ _00253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_95_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11188_ _04918_ mod.u_cpu.rf_ram.memory\[332\]\[0\] _04927_ _04928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_68_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08461__S1 _01838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11736__I _03871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_209_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10139_ _04199_ mod.u_cpu.rf_ram.memory\[497\]\[1\] _04206_ _04208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_67_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_212_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_209_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_209_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09166__I0 mod.u_arbiter.i_wb_cpu_rdt\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14947_ _00801_ net3 mod.u_cpu.rf_ram.memory\[220\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_48_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12768__S _06000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_236_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08669__A2 _02974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13662__A2 _06644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12465__A3 _03377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14878_ _00732_ net3 mod.u_cpu.rf_ram.memory\[248\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_21_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_247_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07341__A2 _01648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_247_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13829_ mod.u_arbiter.i_wb_cpu_rdt\[29\] mod.u_arbiter.i_wb_cpu_rdt\[13\] _06335_
+ _06827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_91_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_250_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07350_ _01657_ _01658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_56_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_206_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_204_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_206_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07281_ _01446_ _01566_ _01588_ _01589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_104_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09876__I _04025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09020_ _03323_ _03324_ _03325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__14723__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_191_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13398__I _06285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09641__I1 mod.u_cpu.rf_ram.memory\[564\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_176_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07396__I _01538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10787__I0 _04637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_176_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_105_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_254_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14873__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09922_ _04057_ _00168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_98_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_258_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__12153__A2 _05568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09853_ _04009_ _00147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_213_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08804_ _01511_ mod.u_cpu.rf_ram.memory\[70\]\[1\] _03110_ _02109_ _03111_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09784_ _03936_ mod.u_cpu.rf_ram.memory\[54\]\[1\] _03955_ _03957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__15229__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08109__A1 _02150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09116__I _03414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07580__A2 _01873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_230_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08735_ _02179_ mod.u_cpu.rf_ram.memory\[252\]\[1\] _03041_ _03042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_3119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13653__A2 _06660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_215_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_199_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08666_ mod.u_cpu.rf_ram.memory\[218\]\[1\] mod.u_cpu.rf_ram.memory\[219\]\[1\] _02294_
+ _02973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_2429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_199_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07999__C _02306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10711__I0 _04593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_214_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_187_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_242_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_199_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14253__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07617_ _01924_ _01925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_54_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_199_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15379__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08597_ _02070_ mod.u_cpu.rf_ram.memory\[260\]\[1\] _02903_ _02904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09609__A1 _03707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13405__A2 _06413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09987__S _04100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_179_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07548_ _01603_ _01856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07479_ mod.u_cpu.raddr\[3\] _01787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_210_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08832__A2 _03131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09786__I _03915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09218_ _03482_ _00037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_167_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_210_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10490_ _04315_ _04443_ _04454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_108_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09149_ mod.u_arbiter.i_wb_cpu_dbus_dat\[3\] _03441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10725__I _04541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13101__I _06017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08596__A1 _01858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12160_ _05588_ _05589_ _05590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_151_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_162_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08691__S1 _02350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11111_ _04862_ mod.u_cpu.rf_ram.memory\[345\]\[1\] _04874_ _04876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_151_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12091_ _05387_ _05543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_162_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14133__S _07053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5000 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13192__I1 mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11042_ _04277_ _04822_ _04828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_5011 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xtiny_user_project_12 io_oeb[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_104_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xtiny_user_project_23 io_oeb[15] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__10155__A1 _04218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_249_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5022 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xtiny_user_project_34 io_oeb[26] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_118_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5033 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_231_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__13892__A2 _06223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5044 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xtiny_user_project_45 io_oeb[37] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_76_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xtiny_user_project_56 io_out[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_5055 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_77_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5066 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xtiny_user_project_67 io_out[23] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_265_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xtiny_user_project_78 io_out[34] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__10950__I0 _04753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtiny_user_project_89 la_data_out[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_5077 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_218_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5088 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14801_ _00655_ net3 mod.u_cpu.rf_ram.memory\[287\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_188_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5099 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_218_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_4376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12993_ _06162_ mod.u_cpu.cpu.genblk3.csr.mcause3_0\[0\] _06164_ _06165_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_3642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14732_ _00586_ net3 mod.u_cpu.rf_ram.memory\[321\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11944_ _05446_ _00801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_79_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13704__C _06320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2930 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10702__I0 _04584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_233_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_205_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08520__A1 _01858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2941 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_206_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2952 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2963 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_232_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_229_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_14663_ _00517_ net3 mod.u_cpu.rf_ram.memory\[356\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11875_ _05396_ _05397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_72_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_221_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2974 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2985 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2996 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14746__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10826_ _04678_ _00451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_13614_ _03313_ _03378_ _06632_ _01285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_14594_ _00448_ net3 mod.u_cpu.rf_ram.memory\[390\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_186_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_207_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_201_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12080__A1 _05535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10757_ _04632_ _00428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_13545_ mod.u_arbiter.i_wb_cpu_dbus_adr\[7\] mod.u_arbiter.i_wb_cpu_dbus_adr\[8\]
+ _06589_ _06591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_201_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08823__A2 _03122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_13476_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[19\] _06538_ _06540_ _03598_ _06544_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__10630__A2 _04528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_185_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10688_ _04579_ mod.u_cpu.rf_ram.memory\[412\]\[1\] _04585_ _04587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08533__C _01683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14896__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15215_ _01068_ net3 mod.u_cpu.rf_ram.memory\[135\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12427_ _05019_ _04442_ _05771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09379__A3 _03586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09623__I1 mod.u_cpu.rf_ram.memory\[566\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12358_ _05724_ _00937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_15146_ _00999_ net3 mod.u_cpu.rf_ram.memory\[161\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_181_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11309_ _04989_ _05011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_15077_ _00931_ net3 mod.u_cpu.rf_ram.memory\[183\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_113_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12289_ _05677_ mod.u_cpu.rf_ram.memory\[18\]\[1\] _05675_ _05678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08339__A1 _02421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07944__I _01827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14028_ _06981_ _06983_ _01348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_68_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09000__A2 mod.u_cpu.cpu.alu.i_rs1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11194__I0 _04918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_214_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_132_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14276__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_255_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_222_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_209_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15521__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08520_ _01858_ _02826_ _02827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_64_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08708__C _02633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08451_ _02630_ _02681_ _02722_ _02757_ _02758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_212_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_251_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07402_ _01509_ _01710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_224_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_260_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08382_ mod.u_cpu.rf_ram.memory\[424\]\[1\] mod.u_cpu.rf_ram.memory\[425\]\[1\] mod.u_cpu.rf_ram.memory\[426\]\[1\]
+ mod.u_cpu.rf_ram.memory\[427\]\[1\] _02688_ _02475_ _02689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__09067__A2 _03369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14060__A2 _06998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_182_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08114__I1 mod.u_cpu.rf_ram.memory\[49\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07333_ _01608_ _01640_ _01641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_52_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14218__S _07106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_177_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09862__I1 mod.u_cpu.rf_ram.memory\[53\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07264_ _01504_ _01572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_164_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09003_ mod.u_cpu.cpu.alu.i_rs1 _03308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_176_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_192_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07195_ _01498_ _01503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_117_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_258_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12374__A2 _03866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_160_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11577__S _05192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07250__A1 _01511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15051__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_259_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_160_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09905_ _04036_ mod.u_cpu.rf_ram.memory\[533\]\[1\] _04042_ _04046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_99_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14619__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13874__A2 _06834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_101_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_219_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09836_ _03945_ _03997_ _03998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_101_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_247_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14123__I0 _07043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09767_ _03944_ _03945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_132_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12201__S _05615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14769__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08718_ _01704_ _03024_ _03025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09698_ _03762_ _03889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_2248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08649_ _02130_ _02955_ _02956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_214_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_70_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_11660_ _05243_ mod.u_cpu.rf_ram.memory\[257\]\[0\] _05247_ _05248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_199_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_230_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10611_ _04255_ _04534_ _04535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11591_ _05194_ mod.u_cpu.rf_ram.memory\[268\]\[1\] _05200_ _05202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_179_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08805__A2 _03108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10999__I0 _04797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_195_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13330_ _06316_ _06426_ _06427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_22_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10542_ _04352_ _04487_ _04488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_155_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_194_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_210_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_183_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13261_ _06126_ mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat\[7\] _06359_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_182_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10473_ _04441_ _00335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_15000_ _00854_ net3 mod.u_cpu.rf_ram.memory\[67\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12212_ mod.u_cpu.rf_ram.memory\[1\]\[1\] _05617_ _05623_ _05625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_157_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11412__I1 _05065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13192_ mod.u_arbiter.i_wb_cpu_rdt\[15\] mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat\[15\]
+ _03499_ _06299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_163_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12143_ _05578_ _00868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_159_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07241__A1 _01505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12670__I _05937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13165__I1 mod.u_cpu.rf_ram.memory\[349\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_235_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12074_ _05521_ mod.u_cpu.rf_ram.memory\[64\]\[0\] _05531_ _05532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_151_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14299__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11286__I _04995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11176__I0 _04918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08416__S1 _02325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15544__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11025_ _04815_ _00513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11876__A1 _05395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10679__A2 _04570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08741__A1 _01978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14114__I0 _07041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_237_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_225_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_206_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_264_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_218_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12976_ _06150_ _06151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_206_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_14715_ _00569_ net3 mod.u_cpu.rf_ram.memory\[330\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_166_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11927_ _05348_ _05434_ _05435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_3494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_178_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_162_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14646_ _00500_ net3 mod.u_cpu.rf_ram.memory\[364\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_127_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11858_ _05384_ _00777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_127_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14042__A2 _06987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_242_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10809_ _04667_ _00445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_11789_ _05329_ mod.u_cpu.rf_ram.memory\[234\]\[1\] _05336_ _05338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_14577_ _00431_ net3 mod.u_cpu.rf_ram.memory\[3\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_159_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13528_ _06580_ _01251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10603__A2 _04528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_201_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08263__C _02469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13459_ _06533_ _01229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__15074__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_138_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15129_ _00982_ net3 mod.u_cpu.rf_ram.memory\[168\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_82_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07951_ _02245_ _02258_ _02259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_142_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13856__A2 _06292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07882_ _02026_ _02190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_214_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_210_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14911__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09621_ _03828_ _03829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_68_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11924__I _05421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10390__I1 mod.u_cpu.rf_ram.memory\[460\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09552_ _03773_ _03774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12667__I0 _05934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08503_ _01520_ _02809_ _02810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_24_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09483_ _01531_ _03708_ _03709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_52_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12292__A1 _05443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07342__C _01615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_197_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_102_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08434_ _02687_ _02733_ _02740_ _01658_ _02741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_212_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_196_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12419__I0 mod.u_cpu.rf_ram.memory\[489\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_212_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_212_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_196_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12044__A1 _05164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08365_ _02026_ _02672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_225_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_211_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07316_ _01556_ mod.u_cpu.rf_ram.memory\[484\]\[0\] _01623_ _01624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_108_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13792__A1 _06425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15417__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08296_ _02066_ _02602_ _02603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_164_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09460__A2 _03337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_178_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07247_ mod.u_cpu.rf_ram.memory\[472\]\[0\] mod.u_cpu.rf_ram.memory\[473\]\[0\] mod.u_cpu.rf_ram.memory\[474\]\[0\]
+ mod.u_cpu.rf_ram.memory\[475\]\[0\] _01540_ _01501_ _01555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_192_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12347__A2 _05703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07178_ _01485_ _01486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_145_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14441__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15567__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08810__I2 mod.u_cpu.rf_ram.memory\[6\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08971__A1 mod.u_cpu.cpu.bufreg2.i_cnt_done vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07774__A2 _02081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11158__I0 _04901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_266_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_232_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14591__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_219_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09819_ _03983_ _00139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_235_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10530__A1 _04439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_246_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12830_ _03781_ _05721_ _06043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2001 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12658__I0 _05923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_185_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2012 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2023 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09304__I _03407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_262_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2034 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_160_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2045 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2056 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12761_ _05997_ _01067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_258_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__11330__I0 _05007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_188_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_265_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2067 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14500_ _00354_ net3 mod.u_cpu.rf_ram.memory\[437\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2078 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11712_ _05254_ _05284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2089 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_215_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15480_ _01252_ net3 mod.u_cpu.rf_ram.memory\[129\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12692_ _04643_ _05952_ _05953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_203_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_199_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_230_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_243_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11643_ _05222_ mod.u_cpu.rf_ram.memory\[25\]\[0\] _05236_ _05237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_187_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14431_ _00285_ net3 mod.u_cpu.rf_ram.memory\[472\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12665__I _05886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13083__I0 _06205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_196_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15097__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_230_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13783__A1 _06739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11574_ _05190_ _00687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_167_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14362_ _00216_ net3 mod.u_cpu.rf_ram.memory\[506\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_195_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13313_ _06338_ _06363_ _06400_ _06410_ _06411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_10525_ _04469_ mod.u_cpu.rf_ram.memory\[438\]\[0\] _04476_ _04477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_14293_ _00147_ net3 mod.u_cpu.rf_ram.memory\[541\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_196_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13244_ _06276_ mod.u_cpu.rf_ram.memory\[93\]\[1\] _06345_ _06347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_109_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10456_ _04176_ _04429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_108_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10349__A1 _04201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07214__A1 _01520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13175_ _06281_ _06282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_124_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10387_ mod.u_cpu.rf_ram.memory\[461\]\[1\] _04383_ _04381_ _04384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07494__I _01752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14934__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12126_ _05566_ mod.u_cpu.rf_ram.memory\[20\]\[1\] _05564_ _05567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07765__A2 _02072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07427__C _01534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13838__A2 _03404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12057_ _05520_ _05521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_96_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11008_ _03931_ _04804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_77_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_226_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_265_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_209_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_179_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12959_ mod.u_arbiter.i_wb_cpu_ibus_adr\[1\] _05783_ _06136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_252_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14314__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07376__S1 _01683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_221_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14015__A2 _06964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14629_ _00483_ net3 mod.u_cpu.rf_ram.memory\[373\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10296__S _04319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_221_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_194_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08274__B _02520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07669__I _01484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_202_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13774__A1 _06289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08150_ mod.u_cpu.rf_ram.memory\[549\]\[0\] _02458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_140_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12577__A2 _05374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_202_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11624__I1 mod.u_cpu.rf_ram.memory\[262\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_187_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14464__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10095__I _03761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08081_ mod.u_cpu.rf_ram.memory\[12\]\[0\] mod.u_cpu.rf_ram.memory\[13\]\[0\] mod.u_cpu.rf_ram.memory\[14\]\[0\]
+ mod.u_cpu.rf_ram.memory\[15\]\[0\] _02266_ _02388_ _02389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__07453__A1 _01759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_220_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13526__A1 _03980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_175_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08721__C _01657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07205__A1 _01511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11001__A2 _04780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_255_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08983_ mod.u_cpu.cpu.branch_op _03254_ _03288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_103_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__10760__A1 _04196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_229_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07934_ _01604_ _02242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_102_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4909 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12888__I0 _06073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07865_ mod.u_cpu.rf_ram.memory\[200\]\[0\] mod.u_cpu.rf_ram.memory\[201\]\[0\] mod.u_cpu.rf_ram.memory\[202\]\[0\]
+ mod.u_cpu.rf_ram.memory\[203\]\[0\] _02171_ _02172_ _02173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_256_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_217_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11560__I0 _05180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08449__B _01591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_228_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09604_ _03802_ mod.u_cpu.rf_ram.memory\[568\]\[0\] _03815_ _03816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_56_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07796_ _01458_ _02104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_83_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_244_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09535_ _03752_ _03758_ _03759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_25_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10115__I1 mod.u_cpu.rf_ram.memory\[500\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_212_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09466_ _03692_ _03693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_262_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__13802__C _06486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_184_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07692__A1 _01711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12017__A1 _05494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08417_ mod.u_cpu.rf_ram.memory\[413\]\[1\] _02724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_240_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14807__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09397_ _03386_ mod.u_scanchain_local.module_data_in\[63\] _03401_ mod.u_arbiter.i_wb_cpu_dbus_adr\[26\]
+ _03634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__13065__I0 _06205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_185_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07579__I _01886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08348_ mod.u_cpu.rf_ram.memory\[494\]\[1\] mod.u_cpu.rf_ram.memory\[495\]\[1\] _01709_
+ _02655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_123_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_193_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08279_ mod.u_cpu.rf_ram.memory\[462\]\[1\] mod.u_cpu.rf_ram.memory\[463\]\[1\] _02585_
+ _02586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_138_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10310_ _04330_ mod.u_cpu.rf_ram.memory\[473\]\[1\] _04328_ _04331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_193_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__14957__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11290_ _04951_ _04999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08619__S1 _02067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11829__I _05328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10241_ _03974_ _04281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_156_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10051__I0 _04140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09992__I0 _04096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10172_ _04232_ _00243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_79_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14980_ _00834_ net3 mod.u_cpu.rf_ram.memory\[60\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12879__I0 _06070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_248_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13931_ _05801_ _06906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_130_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_19_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_235_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_208_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_247_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14337__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13862_ _06814_ _06849_ _06855_ _06704_ _06856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_75_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09034__I mod.u_cpu.cpu.bufreg2.i_cnt_done vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15601_ _01372_ net3 mod.u_cpu.rf_ram.memory\[110\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_263_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12813_ _03774_ _06032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11059__A2 _04704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13793_ _06779_ _06792_ _06793_ _06776_ _06794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_76_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_234_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15532_ _01303_ net3 mod.u_cpu.cpu.immdec.imm30_25\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12744_ _05843_ _05986_ _05987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11854__I1 mod.u_cpu.rf_ram.memory\[6\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13712__C _06135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14487__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08806__C _02677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15463_ _01237_ net3 mod.u_cpu.cpu.ctrl.o_ibus_adr\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07710__C _02005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_179_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12675_ _05934_ mod.u_cpu.rf_ram.memory\[143\]\[0\] _05941_ _05942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_169_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_230_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13756__A1 _01479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14414_ _00268_ net3 mod.u_cpu.rf_ram.memory\[480\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11606__I1 _04954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11626_ _05208_ mod.u_cpu.rf_ram.memory\[262\]\[1\] _05223_ _05225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_169_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15394_ _01169_ net3 mod.u_cpu.rf_ram.memory\[102\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_184_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10034__A3 _03753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14345_ _00199_ net3 mod.u_cpu.rf_ram.memory\[515\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11557_ _05179_ _00681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_239_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10508_ _04453_ mod.u_cpu.rf_ram.memory\[441\]\[0\] _04465_ _04466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_11488_ _05133_ _05131_ _05134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_183_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14276_ _00130_ net3 mod.u_cpu.rf_ram.memory\[54\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_155_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13227_ _03502_ _06334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_10439_ _04418_ _00324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_171_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08113__I _01919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13158_ _06270_ _01191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_124_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_111_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15112__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12109_ _05555_ _00857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13089_ _02287_ _06227_ _06228_ _01164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_266_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_266_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_238_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07650_ _01827_ _01958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_65_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15262__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_207_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07581_ _01849_ _01871_ _01888_ _01889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_230_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_240_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_253_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09320_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[14\] _03569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09112__A1 _03404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13995__A1 mod.u_arbiter.i_wb_cpu_rdt\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_234_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_222_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09251_ _03508_ _03510_ _03511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07620__C _01783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08202_ mod.u_cpu.rf_ram.memory\[565\]\[0\] _02510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_194_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09182_ _03462_ _00020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_193_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_147_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08133_ _02161_ mod.u_cpu.rf_ram.memory\[46\]\[0\] _02440_ _01828_ _02441_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_105_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07426__A1 _01703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_174_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07977__A2 _02284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08064_ _02302_ mod.u_cpu.rf_ram.memory\[76\]\[0\] _02371_ _02372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_174_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07521__S1 _01828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10981__A1 _04784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07285__S0 _01540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_130_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11585__S _05196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_88_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08966_ mod.u_cpu.cpu.immdec.imm11_7\[0\] _03271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_4706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07862__I _01741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15605__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11289__A2 _04997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12486__A1 _05606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07917_ _01518_ _02225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_263_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_217_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08897_ _02471_ _03196_ _03203_ _02518_ _03204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_56_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_257_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09351__A1 _03590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_229_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_217_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07848_ _01635_ _02156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_72_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_245_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_216_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07779_ mod.u_cpu.rf_ram.memory\[180\]\[0\] mod.u_cpu.rf_ram.memory\[181\]\[0\] mod.u_cpu.rf_ram.memory\[182\]\[0\]
+ mod.u_cpu.rf_ram.memory\[183\]\[0\] _02085_ _02086_ _02087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_266_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08537__S0 _01826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09789__I _03960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09518_ _01418_ _01498_ _01518_ _03742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_169_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10790_ _04654_ _00439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_266_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_169_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__07665__A1 _01961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_197_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09449_ _03675_ _03676_ _03677_ _00005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_200_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_200_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_212_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__07760__S1 _02067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12460_ _05792_ _05796_ _05797_ mod.u_arbiter.i_wb_cpu_dbus_dat\[6\] _05798_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_138_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_240_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11411_ _05080_ _00634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_149_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12391_ _03770_ _04142_ _05747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12410__A1 _05759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14136__S _07053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11342_ _04749_ _05011_ _05034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_181_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14130_ _07041_ mod.u_cpu.rf_ram.memory\[118\]\[1\] _07050_ _07052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_138_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_193_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_153_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15135__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_193_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14163__A1 _06062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11273_ _02398_ _04985_ _04986_ _00590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_14061_ _07006_ _07007_ _01357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_181_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_140_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08917__A1 _02471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09029__I _03302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13910__A1 _03679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10224_ _04230_ _04269_ _04270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_13012_ _03837_ _06080_ _06178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09965__I0 _04071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10724__A1 _04184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08393__A2 _02691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10155_ _04218_ _04202_ _04219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15285__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_255_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07772__I _01661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14963_ _00817_ net3 mod.u_cpu.rf_ram.memory\[559\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10086_ _04162_ mod.u_cpu.rf_ram.memory\[504\]\[0\] _04169_ _04170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__13674__B1 _06682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08089__B _02396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13674__C2 _06306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09342__A1 _03568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13914_ _06476_ _06892_ _06893_ _06894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_47_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14894_ _00748_ net3 mod.u_cpu.rf_ram.memory\[237\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_169_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_223_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12229__A1 _05226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13845_ _06775_ _06839_ _06450_ _06840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_222_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_235_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_204_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09699__I _03889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13776_ _06322_ _06714_ _06778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_10988_ _04774_ mod.u_cpu.rf_ram.memory\[363\]\[0\] _04789_ _04790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_200_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_15515_ _01286_ net3 mod.u_cpu.rf_ram.memory\[319\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12727_ _05963_ mod.u_cpu.rf_ram.memory\[78\]\[0\] _05975_ _05976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_95_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_204_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13729__B2 _06735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_175_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15446_ _01220_ net3 mod.u_cpu.cpu.ctrl.o_ibus_adr\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_50_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_12658_ _05923_ mod.u_cpu.rf_ram.memory\[145\]\[1\] _05928_ _05930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_198_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_198_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11609_ _05213_ _00699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_191_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12853__I _06056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15377_ _01152_ net3 mod.u_cpu.rf_ram.memory\[82\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_184_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12589_ _05869_ mod.u_cpu.rf_ram.memory\[156\]\[0\] _05883_ _05884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_172_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14328_ _00182_ net3 mod.u_cpu.rf_ram.memory\[523\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_176_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_117_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11469__I _05118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08271__C _02578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10373__I _04308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_176_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14259_ _00113_ net3 mod.u_cpu.rf_ram.memory\[558\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__14502__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15628__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08908__A1 _02449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13901__A1 _03306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13684__I _06367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_213_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08820_ _02411_ _03126_ _03127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_174_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08751_ _01670_ _03057_ _02230_ _03058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_97_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_245_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_239_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11515__I0 _05147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14652__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07702_ _01581_ _02010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_113_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08682_ _02477_ _02987_ _02988_ _01638_ _02989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_94_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_241_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07633_ _01938_ mod.u_cpu.rf_ram.memory\[310\]\[0\] _01940_ _01783_ _01941_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_80_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_241_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_198_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15008__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13968__A1 mod.u_arbiter.i_wb_cpu_rdt\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07564_ _01851_ _01872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13968__B2 _03444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_179_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09402__I _03637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09303_ _03495_ _03554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_263_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_210_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07495_ mod.u_cpu.rf_ram.memory\[445\]\[0\] _01803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_139_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07111__A3 mod.u_cpu.cpu.csr_d_sel vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07742__S1 _02049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09234_ _03405_ _03495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_194_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15158__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_210_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09165_ _03451_ _03452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__13196__A2 mod.u_arbiter.i_wb_cpu_rdt\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12243__I1 mod.u_cpu.rf_ram.memory\[196\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_222_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08116_ mod.u_cpu.rf_ram.memory\[56\]\[0\] mod.u_cpu.rf_ram.memory\[57\]\[0\] mod.u_cpu.rf_ram.memory\[58\]\[0\]
+ mod.u_cpu.rf_ram.memory\[59\]\[0\] _02242_ _02267_ _02424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_163_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12943__A2 _03458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08998__I1 _03302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09096_ mod.u_cpu.cpu.state.init_done _03391_ _03393_ _03396_ _03397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_107_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08047_ _02135_ mod.u_cpu.rf_ram.memory\[68\]\[0\] _02354_ _02355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_190_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10006__I0 _04096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09947__I0 _04073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11754__I0 _05311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_131_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_5204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07806__B _02113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09998_ _04107_ _04108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_5237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_237_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xtiny_user_project_107 la_data_out[25] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_5259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xtiny_user_project_118 la_data_out[36] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_4514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12459__A1 _03338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xtiny_user_project_129 la_data_out[47] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_08949_ mod.u_cpu.cpu.decode.opcode\[0\] _03254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11506__I0 _05144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_4536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09324__A1 _03436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13120__A2 _04708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09324__B2 mod.u_arbiter.i_wb_cpu_dbus_adr\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11960_ _05457_ _00806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_29_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_151_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10911_ _04172_ _04713_ _04737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_3868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07886__A1 _02191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11891_ _05408_ _05401_ _05409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11682__A2 _05263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_204_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11842__I _05373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_217_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08637__B _02102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13630_ _06485_ _06284_ _06322_ _06305_ _06643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_10842_ _04689_ _00456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_73_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_240_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__12631__A1 _05870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13561_ mod.u_arbiter.i_wb_cpu_dbus_adr\[14\] mod.u_arbiter.i_wb_cpu_dbus_adr\[15\]
+ _06599_ _06600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_198_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10773_ _03895_ _04643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_198_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_160_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15300_ _00060_ net4 mod.u_scanchain_local.module_data_in\[57\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_201_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12512_ _05822_ mod.u_cpu.rf_ram.memory\[168\]\[1\] _05832_ _05834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_12_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13492_ _03624_ _06551_ _06552_ _03631_ _06554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_100_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15231_ _01084_ net3 mod.u_cpu.rf_ram.memory\[229\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_139_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_199_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12443_ _03498_ _05781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_139_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12673__I _05919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08438__I0 mod.u_cpu.rf_ram.memory\[388\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_240_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_199_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09468__B _03694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_201_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11198__A1 _04792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08372__B _02664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10245__I0 _04267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14525__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08063__A1 _02369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15162_ _01015_ net3 mod.u_cpu.rf_ram.memory\[153\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_197_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12374_ _05563_ _03866_ _05736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_165_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_193_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11993__I0 _05470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_176_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_153_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10193__I _03737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14113_ _06903_ _07041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_11325_ _05022_ _05021_ _05023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_153_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07810__A1 _02116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15093_ _00947_ net3 mod.u_cpu.rf_ram.memory\[177\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_101_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11256_ _04973_ _04969_ _04974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_14044_ mod.u_arbiter.i_wb_cpu_dbus_dat\[25\] _06989_ _06995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_140_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__14675__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09563__A1 _03758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10207_ _04245_ mod.u_cpu.rf_ram.memory\[488\]\[1\] _04256_ _04258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_11187_ _04784_ _04926_ _04927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_136_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_121_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10138_ _04207_ _00234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_94_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_227_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_251_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09315__A1 mod.u_arbiter.i_wb_cpu_dbus_adr\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09166__I1 mod.u_arbiter.i_wb_cpu_dbus_dat\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14946_ _00800_ net3 mod.u_cpu.rf_ram.memory\[220\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10069_ _04157_ mod.u_cpu.rf_ram.memory\[507\]\[1\] _04155_ _04158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_209_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11122__A1 _03879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_208_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12465__A4 _05802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_251_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_14877_ _00731_ net3 mod.u_cpu.rf_ram.memory\[253\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_78_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11752__I _03884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_223_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08547__B _01891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13828_ _06283_ _06824_ _06825_ _06642_ _06826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_90_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_204_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07629__A1 _01643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_210_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_13759_ _06492_ _06712_ _06762_ _06475_ _06412_ _06763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_149_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12784__S _06012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15300__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_182_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_149_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07280_ _01536_ _01571_ _01585_ _01587_ _01588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_86_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15429_ _01204_ net3 mod.u_cpu.rf_ram.memory\[95\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09378__B _03616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_191_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08054__A1 _02352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15450__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10936__A1 _04352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14127__A1 _03828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09921_ _04051_ mod.u_cpu.rf_ram.memory\[530\]\[0\] _04056_ _04057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_132_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_217_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13886__B1 _06871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09554__A1 _03775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10831__I _04640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09852_ _03999_ mod.u_cpu.rf_ram.memory\[541\]\[1\] _04007_ _04009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_219_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08803_ _02190_ _03109_ _03110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_252_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09783_ _03956_ _00130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07345__C _01618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08109__A2 _02404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08734_ _02197_ _03040_ _03041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_227_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11113__A1 _04732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08665_ _02561_ _02968_ _02971_ _01696_ _02972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_121_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11662__I _05106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10711__I1 mod.u_cpu.rf_ram.memory\[408\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07616_ _01634_ _01924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_183_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08596_ _01858_ _02902_ _02903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_81_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09132__I mod.u_arbiter.i_wb_cpu_rdt\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_224_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10278__I _04301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07547_ _01854_ _01855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_14_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14548__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08293__A1 _01607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07478_ _01773_ _01777_ _01784_ _01785_ _01786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_195_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_194_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_179_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09217_ mod.u_scanchain_local.module_data_in\[35\] mod.u_arbiter.i_wb_cpu_dbus_dat\[30\]
+ _03479_ _03482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_10_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_259_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__13413__I0 _06351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11103__S _04870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_182_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_148_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09148_ _03440_ _00076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_147_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_194_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_136_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10778__I1 _04532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__14698__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09079_ _03379_ _03304_ _03380_ _03381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_68_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11110_ _04875_ _00538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_151_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12090_ _05542_ _00851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_155_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11041_ _04802_ _04827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_89_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10741__I _04620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5001 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xtiny_user_project_13 io_oeb[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_5012 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10155__A2 _04202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5023 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08899__A3 _03205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtiny_user_project_24 io_oeb[16] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_5034 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xtiny_user_project_35 io_oeb[27] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_103_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xtiny_user_project_46 io_out[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_4300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_77_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5045 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_209_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_190_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07651__S0 _01957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_57 io_out[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_264_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5056 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_162_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5067 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_68 io_out[24] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_58_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5078 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14800_ _00654_ net3 mod.u_cpu.rf_ram.memory\[287\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_4333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xtiny_user_project_79 io_out[35] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__10950__I1 mod.u_cpu.rf_ram.memory\[36\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5089 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12992_ _06163_ _06164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_4366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14731_ _00585_ net3 mod.u_cpu.rf_ram.memory\[322\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_233_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_4399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07859__A1 _02155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11943_ _05426_ mod.u_cpu.rf_ram.memory\[220\]\[1\] _05444_ _05446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_3665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2920 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15323__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2931 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_205_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_260_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08520__A2 _02826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2942 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_205_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14662_ _00516_ net3 mod.u_cpu.rf_ram.memory\[356\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2953 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2964 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11874_ _05386_ _05396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_189_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2975 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2986 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13613_ _03378_ _06631_ _06632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2997 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10825_ _04666_ mod.u_cpu.rf_ram.memory\[38\]\[1\] _04676_ _04678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_186_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14593_ _00447_ net3 mod.u_cpu.rf_ram.memory\[391\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_207_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13801__B1 _06800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_198_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13544_ _06590_ _01257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__15473__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12080__A2 _05471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10756_ _04622_ mod.u_cpu.rf_ram.memory\[400\]\[0\] _04631_ _04632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_71_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_201_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13499__I _06539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_185_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_158_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13475_ _06543_ _01235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_201_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10687_ _04586_ _00404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_127_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15214_ _01067_ net3 mod.u_cpu.rf_ram.memory\[135\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_145_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12426_ _05770_ _00959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_166_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10918__A1 _04741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11966__I0 _05450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_142_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15145_ _00998_ net3 mod.u_cpu.rf_ram.memory\[162\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_126_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12357_ _05711_ mod.u_cpu.rf_ram.memory\[122\]\[1\] _05722_ _05724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_114_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_236_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11308_ _05010_ _00601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_114_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15076_ _00930_ net3 mod.u_cpu.rf_ram.memory\[183\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12288_ _05634_ _05677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_113_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13332__A2 _06326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14027_ mod.u_arbiter.i_wb_cpu_rdt\[19\] _06976_ _06982_ mod.u_arbiter.i_wb_cpu_dbus_dat\[19\]
+ _06983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_136_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_214_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_11239_ _04961_ mod.u_cpu.rf_ram.memory\[324\]\[0\] _04962_ _04963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_141_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_256_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12779__S _06007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_236_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_209_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_209_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14929_ _00783_ net3 mod.u_cpu.rf_ram.memory\[71\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_82_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08277__B _02584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_247_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08450_ _02742_ _02756_ _01483_ _02757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_91_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07401_ _01516_ _01709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08381_ _01879_ _02688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_177_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_211_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07332_ mod.u_cpu.rf_ram.memory\[493\]\[0\] _01640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__09887__I _03995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08275__A1 _01459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_177_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_220_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_32_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_220_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07263_ mod.u_cpu.rf_ram.memory\[464\]\[0\] mod.u_cpu.rf_ram.memory\[465\]\[0\] mod.u_cpu.rf_ram.memory\[466\]\[0\]
+ mod.u_cpu.rf_ram.memory\[467\]\[0\] _01567_ _01570_ _01571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__14840__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09002_ _01430_ _03307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08027__A1 _01693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07194_ mod.u_cpu.rf_ram.memory\[448\]\[0\] mod.u_cpu.rf_ram.memory\[449\]\[0\] mod.u_cpu.rf_ram.memory\[450\]\[0\]
+ mod.u_cpu.rf_ram.memory\[451\]\[0\] _01496_ _01501_ _01502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_192_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07200__I _01507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_191_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_144_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11582__A1 _05110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10385__A2 _04381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14990__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13358__B _06131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11709__I0 _05271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09904_ _02563_ _04042_ _04045_ _00162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__14033__I _06963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_113_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12382__I0 _05729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09127__I mod.u_arbiter.i_wb_cpu_rdt\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09835_ _03991_ _03996_ _03997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_100_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12689__S _05947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15346__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13087__A1 _03941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09766_ _03697_ _03944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13805__C _06776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_262_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_215_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08717_ mod.u_cpu.rf_ram.memory\[231\]\[1\] _03024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_2205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_265_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_215_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09697_ _03888_ _00112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_55_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_242_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14370__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_2249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10696__I0 _04584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08648_ mod.u_cpu.rf_ram.memory\[165\]\[1\] _02955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_1515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_54_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__15496__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_26_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_203_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_199_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13821__B _06332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08579_ _01711_ _02885_ _02886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10937__S _04754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_23_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_211_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10610_ _04436_ _04534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08266__A1 _02472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11590_ _05201_ _00692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_195_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_167_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10541_ _04442_ _04487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_167_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_202_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13260_ _06357_ _06358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_108_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10472_ _04430_ mod.u_cpu.rf_ram.memory\[447\]\[1\] _04438_ _04441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_157_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12211_ _05624_ _00890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_203_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_194_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13191_ _05782_ _03456_ _06297_ _06298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_136_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_191_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08650__B _02956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_237_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12142_ _05575_ mod.u_cpu.rf_ram.memory\[75\]\[0\] _05577_ _05578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_194_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_237_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13268__B _06365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09518__A1 _01418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12073_ _05417_ _05388_ _05531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11325__A1 _05022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_249_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11024_ _04797_ mod.u_cpu.rf_ram.memory\[358\]\[1\] _04813_ _04815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_1_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11876__A2 _05397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_265_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14114__I1 mod.u_cpu.rf_ram.memory\[87\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_49_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14713__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12825__A1 _03770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12975_ _03389_ mod.u_cpu.cpu.state.o_cnt\[2\] _06150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_4196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_206_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_233_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_14714_ _00568_ net3 mod.u_cpu.rf_ram.memory\[330\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_261_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_206_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11926_ _04994_ _05433_ _05434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_3484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_244_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14645_ _00499_ net3 mod.u_cpu.rf_ram.memory\[365\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14863__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11857_ _05383_ mod.u_cpu.rf_ram.memory\[6\]\[1\] _05381_ _05384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_2794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_221_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_92_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_220_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08257__A1 _02527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10808_ _04666_ mod.u_cpu.rf_ram.memory\[392\]\[1\] _04664_ _04667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_14576_ _00430_ net3 mod.u_cpu.rf_ram.memory\[3\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_159_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11788_ _05337_ _00754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_198_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_203_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09500__I _03725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08544__C _01492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13527_ _06578_ mod.u_cpu.rf_ram.memory\[129\]\[0\] _06579_ _06580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_10739_ _04619_ _00423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_174_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15219__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13458_ _03552_ _06531_ _06532_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[13\] _06533_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_220_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11678__S _05259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12409_ _05487_ _05759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_126_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12861__I _03338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10582__S _04512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13389_ _06377_ _03449_ _06484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_138_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11564__A1 _04766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15128_ _00981_ net3 mod.u_cpu.rf_ram.memory\[168\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_173_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14243__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11477__I _05124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15369__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10381__I _04378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07950_ mod.u_cpu.rf_ram.memory\[245\]\[0\] _02258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_15059_ _00913_ net3 mod.u_cpu.rf_ram.memory\[190\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_99_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11316__A1 _04732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07881_ mod.u_cpu.rf_ram.memory\[222\]\[0\] mod.u_cpu.rf_ram.memory\[223\]\[0\] _02048_
+ _02189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_229_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_228_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09620_ _03827_ _03828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_56_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14393__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13069__A1 _05742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_255_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07690__I _01752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_244_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08719__C _02154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09551_ _03695_ _03773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07623__C _01812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12667__I1 mod.u_cpu.rf_ram.memory\[121\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08502_ mod.u_cpu.rf_ram.memory\[325\]\[1\] _02809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_224_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12101__I _05549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09482_ _01659_ _03703_ _03708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12292__A2 _05668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_212_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_251_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08433_ _02654_ _02736_ _02739_ _02730_ _02740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_197_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12419__I1 _05765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08364_ _02638_ mod.u_cpu.rf_ram.memory\[484\]\[1\] _02670_ _02671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__13241__A1 _03771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_177_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_177_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_149_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10055__A1 _04013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_177_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09996__A1 _03702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07315_ _01573_ _01622_ _01623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_165_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10556__I _04496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_221_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08295_ mod.u_cpu.rf_ram.memory\[455\]\[1\] _02602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_192_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07246_ _01489_ _01535_ _01553_ _01554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_118_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07177_ _01484_ _01485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_145_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_219_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_160_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__14736__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12355__I0 _05713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_247_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09818_ mod.u_cpu.rf_ram.memory\[545\]\[1\] _03929_ _03981_ _03983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09920__A1 _03859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12807__A1 _05948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09749_ mod.u_cpu.rf_ram.memory\[553\]\[1\] _03929_ _03926_ _03930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_41_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14886__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_228_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__13855__I0 mod.u_arbiter.i_wb_cpu_rdt\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2002 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2013 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2024 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_243_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_215_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08487__A1 _01496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2035 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12760_ _05992_ mod.u_cpu.rf_ram.memory\[135\]\[0\] _05996_ _05997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_215_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2046 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2057 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11330__I1 mod.u_cpu.rf_ram.memory\[310\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2068 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11711_ _03803_ _05283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2079 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12691_ _03723_ _05319_ _05952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_230_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_203_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08645__B _02951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14430_ _00284_ net3 mod.u_cpu.rf_ram.memory\[472\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_202_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11642_ _05110_ _04026_ _05236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_243_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_230_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13783__A2 mod.u_arbiter.i_wb_cpu_rdt\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14361_ _00215_ net3 mod.u_cpu.rf_ram.memory\[507\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10466__I _04435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11573_ _05178_ mod.u_cpu.rf_ram.memory\[271\]\[1\] _05188_ _05190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_204_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_183_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_211_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13312_ _06401_ _06408_ _06409_ _06410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__12991__B1 _03337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10524_ _04180_ _04464_ _04476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_182_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14292_ _00146_ net3 mod.u_cpu.rf_ram.memory\[541\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__14266__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_171_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13243_ _06346_ _01200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__15511__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_196_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10455_ _04428_ _00330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_183_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11546__A1 _05037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07775__I _01785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13174_ mod.u_arbiter.i_wb_cpu_rdt\[10\] mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat\[10\]
+ _05781_ _06281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_124_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07214__A2 _01521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08411__A1 _02656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07845__S0 _02151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10386_ _03928_ _04383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_12125_ _05549_ _05566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_96_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_250_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12056_ _05309_ _05520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_172_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_81_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_266_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11007_ _04802_ _04803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_78_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_266_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_266_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_237_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_226_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_93_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_206_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11961__S _05456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_248_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08478__A1 _01875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_12958_ _06134_ _06135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_234_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_233_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_206_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11909_ _04300_ _05371_ _05421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_2580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12889_ _06082_ _01110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15041__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14628_ _00482_ net3 mod.u_cpu.rf_ram.memory\[373\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_61_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_221_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09230__I mod.u_arbiter.i_wb_cpu_ibus_adr\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14609__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11085__I0 _04841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14559_ _00413_ net3 mod.u_cpu.rf_ram.memory\[408\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_174_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08080_ _02126_ _02388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10832__I0 _04682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08650__A1 _02129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_228_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15191__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13526__A2 _05373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11537__A1 _01982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07685__I _01645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14759__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12585__I0 _05874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07205__A2 _01512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08402__A1 _02654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08982_ mod.u_cpu.cpu.decode.co_mem_word mod.u_cpu.cpu.csr_d_sel _03287_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__10760__A2 _03969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09606__S _03815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07933_ _02170_ _02233_ _02240_ _02168_ _02241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_130_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_229_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_1243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07864_ _01614_ _02172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_56_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09603_ _03814_ _03805_ _03815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07795_ _02089_ _02101_ _02102_ _02103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_84_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_225_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09534_ _03757_ _03758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_43_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08469__A1 _01852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_225_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09465_ _03292_ _03692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_149_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_212_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_212_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_184_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08416_ mod.u_cpu.rf_ram.memory\[408\]\[1\] mod.u_cpu.rf_ram.memory\[409\]\[1\] mod.u_cpu.rf_ram.memory\[410\]\[1\]
+ mod.u_cpu.rf_ram.memory\[411\]\[1\] _02225_ _02325_ _02723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__12017__A2 _05471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_200_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09396_ _03631_ _03627_ _03493_ _03633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__14289__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_225_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08184__C _02491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15534__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08347_ _02218_ _02654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_149_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10823__I0 _04663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08641__A1 _02111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08278_ _01636_ _02585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_138_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07229_ _01515_ _01537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_138_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11528__A1 _04741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_180_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_164_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11111__S _04874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10240_ _04280_ _00263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_65_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10171_ mod.u_cpu.rf_ram.memory\[493\]\[1\] _04111_ _04229_ _04232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_78_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09992__I1 mod.u_cpu.rf_ram.memory\[518\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_191_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_266_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_191_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_232_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__12450__B _05787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13930_ _06905_ _01328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_219_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_208_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11700__A1 _04859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13861_ _06853_ _06854_ _06855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_35_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15600_ _01371_ net3 mod.u_cpu.rf_ram.memory\[110\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_216_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12812_ _04844_ _06030_ _06031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_262_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15064__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08004__S0 _02294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13792_ _06425_ _06373_ _06402_ _06683_ _06793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_90_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_215_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12500__I0 _05822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_216_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15531_ _01302_ net3 mod.u_cpu.cpu.immdec.imm30_25\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12743_ _03790_ _05552_ _05986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_203_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07132__A1 _01439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_231_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15462_ _01236_ net3 mod.u_cpu.cpu.ctrl.o_ibus_adr\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_203_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12674_ _04913_ _05940_ _05941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09050__I _03250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_179_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08094__C _02185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14413_ _00267_ net3 mod.u_cpu.rf_ram.memory\[481\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11625_ _05224_ _00704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_187_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13756__A2 _06657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15393_ _01168_ net3 mod.u_cpu.rf_ram.memory\[102\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_196_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11767__A1 _05322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_204_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14344_ _00198_ net3 mod.u_cpu.rf_ram.memory\[515\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__14901__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11556_ _05178_ mod.u_cpu.rf_ram.memory\[274\]\[1\] _05175_ _05179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_128_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08822__C _02415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10507_ _04163_ _04464_ _04465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13508__A2 _03325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_195_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10924__I _04541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14275_ _00129_ net3 mod.u_cpu.rf_ram.memory\[550\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11487_ _05132_ _05133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13300__I _06397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13226_ _06139_ _06332_ _06333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_109_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10438_ _04400_ mod.u_cpu.rf_ram.memory\[452\]\[0\] _04417_ _04418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_87_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12192__A1 _05334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13157_ mod.u_arbiter.i_wb_cpu_rdt\[29\] mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat\[13\]
+ _06268_ _06270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10369_ _04311_ _04370_ _04371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12108_ _05550_ mod.u_cpu.rf_ram.memory\[211\]\[1\] _05553_ _05555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_69_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13088_ _06032_ _06227_ _06228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_215_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12039_ _05443_ _03810_ _05509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08699__A1 _02190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15407__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_226_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_265_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_254_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07580_ _01872_ _01873_ _01885_ _01887_ _01888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_19_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13444__B2 mod.u_cpu.cpu.ctrl.o_ibus_adr\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09112__A2 _03408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_222_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14431__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__13995__A2 _06952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15557__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09250_ _03509_ _03510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_34_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08201_ _01682_ _02509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09181_ mod.u_arbiter.i_wb_cpu_rdt\[17\] mod.u_arbiter.i_wb_cpu_dbus_dat\[14\] _03459_
+ _03462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_159_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_194_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_222_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11758__A1 _05187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_187_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_239_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08132_ _01819_ _02439_ _02440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_146_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14581__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10805__I0 _04663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_175_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15549__D _01320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_174_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_179_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08063_ _02369_ _02370_ _02371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_147_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10981__A2 _04759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08304__I _02350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_255_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07729__A3 _02036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_216_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_192_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07285__S1 _01570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_170_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_88_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13366__B _06330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08965_ _03269_ mod.u_cpu.cpu.state.o_cnt\[2\] _03270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_233_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_4707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07916_ _01651_ _02223_ _02224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__14041__I _06970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15087__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08896_ _02476_ _03199_ _03202_ _02489_ _03203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_111_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12486__A2 _05767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_256_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07847_ _02154_ _02155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_17_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_244_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_84_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08974__I mod.u_cpu.cpu.bufreg.lsb\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12238__A2 _05641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07778_ _01854_ _02086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_37_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09517_ _01461_ _01778_ _03741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__08907__C _02467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08537__S1 _02164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07811__C _01771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07114__A1 _01421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_262_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_213_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11997__A1 _05019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09448_ _03334_ _03668_ _03677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__14924__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_240_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_149_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09379_ _03602_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[20\] _03586_ _03594_ _03618_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__10945__S _04760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11410_ mod.u_cpu.rf_ram.memory\[297\]\[0\] _04954_ _05079_ _05080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12797__I0 _06010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12390_ _05746_ _00947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_166_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12410__A2 _05758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_193_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11341_ _05033_ _00611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_193_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07539__B _01485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14060_ mod.u_arbiter.i_wb_cpu_rdt\[28\] _06998_ _07004_ mod.u_arbiter.i_wb_cpu_dbus_dat\[28\]
+ _07007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_180_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11272_ _04746_ _04985_ _04986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_152_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14163__A2 _06568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_180_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07258__C _01552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13371__B1 _06465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13011_ _06177_ _01137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_134_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08917__A2 _03216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10223_ _04108_ _04228_ _04269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_106_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14304__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10724__A2 _04574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10154_ _03885_ _04218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_95_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11575__I _05119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_248_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14962_ _00816_ net3 mod.u_cpu.rf_ram.memory\[559\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_66_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13674__A1 _06304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10085_ _04168_ _04164_ _04169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13674__B2 _06661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13913_ _06398_ _06452_ _06695_ _06893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_130_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14454__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_247_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14893_ _00747_ net3 mod.u_cpu.rf_ram.memory\[239\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_130_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_236_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_210_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13844_ _06367_ _06743_ _06839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_74_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_263_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12229__A2 _05594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13775_ _06776_ _06777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_10987_ _04238_ _04788_ _04789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11988__A1 _05448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11016__S _04809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_204_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12726_ _03885_ _05576_ _05975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_15514_ _01285_ net3 mod.u_cpu.cpu.alu.cmp_r vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08853__A1 _01608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_245_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_231_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15445_ _01219_ net3 mod.u_cpu.cpu.ctrl.o_ibus_adr\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_230_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12657_ _05929_ _01031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_188_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11608_ mod.u_cpu.rf_ram.memory\[265\]\[1\] _05065_ _05211_ _05213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08605__A1 _01738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15376_ _01151_ net3 mod.u_cpu.rf_ram.memory\[79\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_128_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09653__I0 _03832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12588_ _05443_ _05882_ _05883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_117_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11460__I0 _05108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14327_ _00181_ net3 mod.u_cpu.rf_ram.memory\[524\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11539_ _05167_ _00675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_128_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14258_ _00112_ net3 mod.u_cpu.rf_ram.memory\[558\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_171_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13209_ _06117_ _06300_ _06316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08908__A2 _03207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13901__A2 _06881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14189_ _07090_ _01402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_174_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_252_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11912__A1 _04845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07592__A1 _01874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08750_ mod.u_cpu.rf_ram.memory\[104\]\[1\] mod.u_cpu.rf_ram.memory\[105\]\[1\] mod.u_cpu.rf_ram.memory\[106\]\[1\]
+ mod.u_cpu.rf_ram.memory\[107\]\[1\] _02106_ _02107_ _03057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_26_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08216__S0 _02494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13665__A1 _06338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_238_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_266_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07701_ _01978_ _01990_ _02008_ _02009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_113_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_266_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08681_ _02632_ mod.u_cpu.rf_ram.memory\[208\]\[1\] _02988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_65_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_226_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07632_ _01507_ _01939_ _01940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_81_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13417__A1 _05732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14947__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_253_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__13968__A2 _06938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07563_ _01852_ _01853_ _01869_ _01870_ _01871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__14090__A1 _07026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_263_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09302_ _03552_ _03549_ _03553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_62_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_250_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_210_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07494_ _01752_ _01802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__08844__A1 _02578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_222_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07203__I _01510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09892__I0 _04036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_179_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09233_ _03491_ _03494_ _00040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_167_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12779__I0 _05998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09164_ _03413_ _03451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_182_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08115_ mod.u_cpu.rf_ram.memory\[60\]\[0\] mod.u_cpu.rf_ram.memory\[61\]\[0\] mod.u_cpu.rf_ram.memory\[62\]\[0\]
+ mod.u_cpu.rf_ram.memory\[63\]\[0\] _02369_ _02218_ _02423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_175_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__14036__I _06914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_175_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09095_ _03394_ _03395_ _03396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_174_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14327__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_190_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08046_ _02266_ _02353_ _02354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_190_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09021__A1 _03298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11754__I1 mod.u_cpu.rf_ram.memory\[238\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_192_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_5205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__14477__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09997_ _04106_ _04107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_131_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_95_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xtiny_user_project_108 la_data_out[26] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_4504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08948_ _01422_ _03253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_4515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xtiny_user_project_119 la_data_out[37] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__12459__A2 _03668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_257_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_229_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08879_ _03176_ _03185_ _02609_ _03186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_3825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08918__B _01447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_229_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10910_ _04736_ _00477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_245_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07886__A2 _02192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11890_ _03973_ _05408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_151_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10841_ _04679_ mod.u_cpu.rf_ram.memory\[386\]\[0\] _04688_ _04689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_60_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_13560_ _06583_ _06599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_164_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10772_ _04642_ _00433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_201_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12631__A2 _03886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09883__I0 _04023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_201_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07113__I mod.u_cpu.cpu.branch_op vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07194__S0 _01496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_241_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_198_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12511_ _05833_ _00981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_9_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11690__I0 _05268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_212_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10493__I1 mod.u_cpu.rf_ram.memory\[444\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15102__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_233_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13491_ _06553_ _01241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_15230_ _01083_ net3 mod.u_cpu.rf_ram.memory\[229\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_40_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12442_ _01433_ _05780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_173_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09635__I0 _03832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_200_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08372__C _02678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15161_ _01014_ net3 mod.u_cpu.rf_ram.memory\[154\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10474__I _04435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_197_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12373_ _05735_ _00941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12934__A3 mod.timer_irq vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15252__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14112_ _07040_ _01375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_11324_ _04541_ _05022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_126_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15092_ _00946_ net3 mod.u_cpu.rf_ram.memory\[177\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_180_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14043_ _06992_ _06994_ _01352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_113_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11255_ _04125_ _04973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_140_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_153_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07783__I _01671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10206_ _04257_ _00252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09563__A2 _03782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11186_ _04905_ _04926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_122_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10137_ _04193_ mod.u_cpu.rf_ram.memory\[497\]\[0\] _04206_ _04207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_209_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_209_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09315__A2 _03564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_236_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14945_ _00799_ net3 mod.u_cpu.rf_ram.memory\[169\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10068_ _04090_ _04157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_47_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_209_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12170__I1 _05468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_208_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14876_ _00730_ net3 mod.u_cpu.rf_ram.memory\[253\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_91_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_235_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_217_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10881__A1 _04315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13827_ _06319_ _06324_ _06643_ _06825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_1_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14072__A1 _03858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_232_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_206_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07629__A2 mod.u_cpu.rf_ram.memory\[308\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08826__A1 _02406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13758_ mod.u_arbiter.i_wb_cpu_rdt\[19\] mod.u_arbiter.i_wb_cpu_rdt\[3\] _03509_
+ _06762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_189_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_204_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_204_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12709_ _05870_ _04668_ _05964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_231_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13689_ _06695_ _06698_ _06699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_143_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15428_ _01203_ net3 mod.u_cpu.rf_ram.memory\[92\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09626__I0 _03832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_191_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08282__C _02188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15359_ _01134_ net3 mod.u_cpu.cpu.genblk3.csr.mcause3_0\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08054__A2 _02355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_176_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14127__A2 _05631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_236_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13695__I _05787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_176_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09920_ _03859_ _04038_ _04056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_116_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_256_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13886__A1 _06382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09851_ _02573_ _04007_ _04008_ _00146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_59_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08802_ mod.u_cpu.rf_ram.memory\[71\]\[1\] _03109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_150_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12104__I _05432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09782_ _03916_ mod.u_cpu.rf_ram.memory\[54\]\[0\] _03955_ _03956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_258_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_239_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08733_ mod.u_cpu.rf_ram.memory\[253\]\[1\] _03040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_22_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_230_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12161__I1 _05437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12040__S _05509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08664_ _02566_ mod.u_cpu.rf_ram.memory\[222\]\[1\] _02970_ _01703_ _02971_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_26_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_241_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_215_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07615_ _01643_ mod.u_cpu.rf_ram.memory\[316\]\[0\] _01922_ _01923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_148_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_198_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15125__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_214_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08595_ mod.u_cpu.rf_ram.memory\[261\]\[1\] _02902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__14063__A1 mod.u_arbiter.i_wb_cpu_rdt\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08117__I0 _02420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08029__I _02057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07546_ _01499_ _01854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08817__A1 _02369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_222_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09490__A1 _03664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07477_ _01765_ _01785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_139_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15275__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09216_ _03481_ _00036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_167_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_210_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09617__I0 _03800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_182_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09147_ mod.u_arbiter.i_wb_cpu_rdt\[5\] _03438_ _03439_ _03440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_148_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13819__B _06779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09078_ mod.u_cpu.cpu.alu.add_cy_r _03356_ _03380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_151_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12129__A1 _05300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_190_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13177__I0 mod.u_arbiter.i_wb_cpu_rdt\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08029_ _02057_ _02337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_122_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13877__A1 mod.u_cpu.cpu.immdec.imm24_20\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11040_ _04826_ _00517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_5002 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xtiny_user_project_14 io_oeb[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_5013 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xtiny_user_project_25 io_oeb[17] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_5024 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_118_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_36 io_oeb[28] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_5035 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_49_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5046 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_130_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_47 io_out[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_58 io_out[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_5057 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07651__S1 _01958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_218_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xtiny_user_project_69 io_out[25] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_40_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5068 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_162_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5079 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12991_ _06062_ _03375_ _03337_ _03336_ _06163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XTAP_4356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07308__A1 _01577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14730_ _00584_ net3 mod.u_cpu.rf_ram.memory\[322\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11942_ _05445_ _00800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_73_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2910 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_3666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2921 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_206_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2932 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_217_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14661_ _00515_ net3 mod.u_cpu.rf_ram.memory\[357\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2943 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10469__I _04043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10863__A1 _04700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11873_ _03940_ _05395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_2954 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14054__A1 _07001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2965 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_221_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2976 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13612_ _06624_ _06628_ _06629_ _06630_ _06631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_214_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2987 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10824_ _04677_ _00450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__15618__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08808__A1 _02337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2998 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14592_ _00446_ net3 mod.u_cpu.rf_ram.memory\[391\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_60_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_260_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13801__B2 _06801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_213_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_201_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13543_ mod.u_arbiter.i_wb_cpu_dbus_adr\[6\] mod.u_arbiter.i_wb_cpu_dbus_adr\[7\]
+ _06589_ _06590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_201_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09479__B _01440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10755_ _04209_ _04623_ _04631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_203_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08383__B _02077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_199_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13474_ _03588_ _06538_ _06540_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[19\] _06543_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_199_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10686_ _04584_ mod.u_cpu.rf_ram.memory\[412\]\[0\] _04585_ _04586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_127_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15213_ _01066_ net3 mod.u_cpu.rf_ram.memory\[80\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_199_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__11415__I0 _05071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14642__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12425_ _05761_ mod.u_cpu.rf_ram.memory\[174\]\[1\] _05768_ _05770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_12_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15144_ _00997_ net3 mod.u_cpu.rf_ram.memory\[162\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_126_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12356_ _05723_ _00936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_153_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13317__B1 _06411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13168__I0 _06276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11307_ _04999_ mod.u_cpu.rf_ram.memory\[314\]\[1\] _05008_ _05010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08830__C _01830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15075_ _00929_ net3 mod.u_cpu.rf_ram.memory\[184\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_181_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12287_ _05676_ _00914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_141_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14792__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14026_ _06970_ _06982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_113_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_206_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11238_ _04821_ _04945_ _04962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_253_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11964__S _05459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11169_ _04901_ mod.u_cpu.rf_ram.memory\[335\]\[0\] _04914_ _04915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_110_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_228_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_209_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15148__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11763__I _05252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_36_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14928_ _00782_ net3 mod.u_cpu.rf_ram.memory\[71\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_48_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_264_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_110_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_236_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_223_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14859_ _00713_ net3 mod.u_cpu.rf_ram.memory\[24\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__14045__A1 mod.u_arbiter.i_wb_cpu_rdt\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14045__B2 mod.u_arbiter.i_wb_cpu_dbus_dat\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07400_ _01705_ mod.u_cpu.rf_ram.memory\[412\]\[0\] _01707_ _01708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__15298__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08380_ _02591_ _02687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_91_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09847__I0 _03999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_189_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_205_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_220_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07331_ mod.u_cpu.rf_ram.memory\[488\]\[0\] mod.u_cpu.rf_ram.memory\[489\]\[0\] mod.u_cpu.rf_ram.memory\[490\]\[0\]
+ mod.u_cpu.rf_ram.memory\[491\]\[0\] _01636_ _01638_ _01639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__12594__I _05886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08114__I3 mod.u_cpu.rf_ram.memory\[51\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_260_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_143_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07262_ _01569_ _01570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_192_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09001_ _03299_ _03306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_192_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11406__I0 _05069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_145_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08027__A2 _02322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07193_ _01500_ _01501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_145_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_247_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13159__I0 mod.u_arbiter.i_wb_cpu_rdt\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11582__A2 _03797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08740__C _01870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12035__S _05506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13859__B2 _06464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12906__I0 _06088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09903_ _04044_ _04042_ _04045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_116_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_59_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12531__A1 _05593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09834_ _03995_ _03996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_115_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10393__I0 _04387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09765_ _03834_ _03942_ _03943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_74_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_230_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08716_ _01608_ mod.u_cpu.rf_ram.memory\[228\]\[1\] _03022_ _03023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_132_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09696_ _03877_ mod.u_cpu.rf_ram.memory\[558\]\[0\] _03887_ _03888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10145__I0 _04199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14515__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_2239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10845__A1 _04285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08647_ mod.u_cpu.rf_ram.memory\[160\]\[1\] mod.u_cpu.rf_ram.memory\[161\]\[1\] mod.u_cpu.rf_ram.memory\[162\]\[1\]
+ mod.u_cpu.rf_ram.memory\[163\]\[1\] _02125_ _02127_ _02954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_254_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_199_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07710__A1 _01961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_215_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_215_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_203_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_82_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_81_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08578_ mod.u_cpu.rf_ram.memory\[285\]\[1\] _02885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_39_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_242_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_148_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08915__C _02515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__11645__I0 _05234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_223_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07529_ _01510_ _01837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__14665__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_195_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_211_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__11114__S _04877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_210_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10540_ _04452_ _04486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_128_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_211_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_241_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_157_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_196_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10471_ _01808_ _04438_ _04440_ _00334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_109_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12210_ mod.u_cpu.rf_ram.memory\[1\]\[0\] _05622_ _05623_ _05624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_136_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13190_ _06116_ mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat\[14\] _06297_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_136_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12770__A1 _04955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12141_ _04930_ _05576_ _05577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_191_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_150_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12072_ _05530_ _00845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_89_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11325__A2 _05021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11023_ _04814_ _00512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13570__I0 mod.u_arbiter.i_wb_cpu_dbus_adr\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_264_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12974_ _06149_ _01128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_252_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15440__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_218_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_205_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14713_ _00567_ net3 mod.u_cpu.rf_ram.memory\[331\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__14027__A1 mod.u_arbiter.i_wb_cpu_rdt\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11925_ _05432_ _05433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07701__A1 _01978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11856_ _05328_ _05383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_14644_ _00498_ net3 mod.u_cpu.rf_ram.memory\[365\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_82_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_207_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10807_ _04640_ _04666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_14575_ _00429_ net3 mod.u_cpu.rf_ram.memory\[400\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11787_ _05311_ mod.u_cpu.rf_ram.memory\[234\]\[0\] _05336_ _05337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_202_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08257__A2 mod.u_cpu.rf_ram.memory\[532\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15590__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_201_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10738_ _04608_ mod.u_cpu.rf_ram.memory\[403\]\[1\] _04617_ _04619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_13526_ _03980_ _05373_ _06579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_185_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_242_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11959__S _05456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13457_ _06513_ _06532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_127_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10669_ _04573_ _00399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_127_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12408_ _05187_ _05757_ _05758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12061__I0 _05518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13388_ _06482_ _06483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_127_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_177_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07768__A1 _02074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15127_ _00980_ net3 mod.u_cpu.rf_ram.memory\[16\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_154_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12339_ _05711_ mod.u_cpu.rf_ram.memory\[183\]\[1\] _05707_ _05712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_126_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15058_ _00912_ net3 mod.u_cpu.rf_ram.memory\[190\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08980__A3 mod.u_cpu.cpu.genblk3.csr.o_new_irq vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_214_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13973__I _06914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14009_ mod.u_arbiter.i_wb_cpu_dbus_dat\[16\] _06966_ _06969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13561__I0 mod.u_arbiter.i_wb_cpu_dbus_adr\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_256_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07880_ _01582_ _02188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08812__S0 _02266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10375__I0 _04365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14538__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13069__A2 _06193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_249_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07940__A1 _02244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07791__I1 mod.u_cpu.rf_ram.memory\[189\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09550_ _03767_ _03771_ _03772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10127__I0 _04199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_209_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08501_ mod.u_cpu.rf_ram.memory\[320\]\[1\] mod.u_cpu.rf_ram.memory\[321\]\[1\] mod.u_cpu.rf_ram.memory\[322\]\[1\]
+ mod.u_cpu.rf_ram.memory\[323\]\[1\] _01920_ _02666_ _02808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_236_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__14688__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09481_ mod.u_cpu.cpu.immdec.imm11_7\[0\] _01441_ _03706_ _03707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_58_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_224_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08432_ _02692_ mod.u_cpu.rf_ram.memory\[406\]\[1\] _02738_ _01918_ _02739_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_91_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_212_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_211_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_168_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08363_ _01561_ _02669_ _02670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09445__A1 _01451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13213__I _06118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07314_ mod.u_cpu.rf_ram.memory\[485\]\[0\] _01622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_108_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_260_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10055__A2 _03859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08294_ _02585_ mod.u_cpu.rf_ram.memory\[452\]\[1\] _02600_ _02601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_220_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07245_ _01536_ _01541_ _01549_ _01552_ _01553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_165_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_192_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08751__B _02230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_178_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_191_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_164_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_180_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07176_ _01450_ _01456_ _01484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_106_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11668__I _05253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08470__C _01849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_195_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_258_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08042__I _01637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__12355__I1 mod.u_cpu.rf_ram.memory\[122\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08184__A1 _02471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15463__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09817_ _03982_ _00138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09920__A2 _04038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07931__A1 _02179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_262_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_189_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11109__S _04874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_234_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09748_ _03928_ _03929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_189_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12807__A2 _06027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13855__I1 mod.u_arbiter.i_wb_cpu_rdt\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2003 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2014 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_261_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11866__I0 _05383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13832__B _03679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2025 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09679_ _03847_ mod.u_cpu.rf_ram.memory\[560\]\[0\] _03874_ _03875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__14009__A1 mod.u_arbiter.i_wb_cpu_dbus_dat\[16\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2036 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08487__A2 mod.u_cpu.rf_ram.memory\[358\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2047 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_215_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11710_ _05282_ _00731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_55_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2058 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2069 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_226_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12690_ _05951_ _01042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12448__B _05785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08645__C _02141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11641_ _05235_ _00709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10747__I _04578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09436__A1 mod.u_cpu.cpu.state.init_done vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_204_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_196_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14360_ _00214_ net3 mod.u_cpu.rf_ram.memory\[507\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11572_ _02028_ _05188_ _05189_ _00686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_168_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08217__I _02454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_168_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07121__I mod.u_cpu.cpu.csr_d_sel vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13311_ _06134_ _06409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_10523_ _04475_ _00351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12991__A1 _06062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14291_ _00145_ net3 mod.u_cpu.rf_ram.memory\[542\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_155_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13242_ _06273_ mod.u_cpu.rf_ram.memory\[93\]\[0\] _06345_ _06346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_143_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10454_ _04423_ mod.u_cpu.rf_ram.memory\[44\]\[0\] _04427_ _04428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_136_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12743__A1 _03790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_182_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13173_ mod.u_cpu.cpu.bufreg.i_sh_signed _06140_ _06280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_237_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08411__A2 mod.u_cpu.rf_ram.memory\[446\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10385_ _01542_ _04381_ _04382_ _00306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07845__S1 _02152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12124_ _05565_ _00862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_97_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_238_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12055_ _05519_ _00839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_137_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_265_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11006_ _04620_ _04802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_42_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09372__B1 _03517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_266_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07724__C _02005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_266_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14830__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_253_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09712__S _03897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_218_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11857__I0 _05383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08478__A2 mod.u_cpu.rf_ram.memory\[366\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12957_ _06064_ _06133_ _06134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_3271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09675__A1 _03870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_234_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11908_ _05420_ _00791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_34_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14980__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12888_ _06073_ mod.u_cpu.rf_ram.memory\[89\]\[0\] _06081_ _06082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_2592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13759__B1 _06762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14627_ _00481_ net3 mod.u_cpu.rf_ram.memory\[374\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11839_ _03662_ _04223_ _03753_ _05371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10037__A2 _04132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_193_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_159_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14558_ _00412_ net3 mod.u_cpu.rf_ram.memory\[408\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_159_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15336__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13509_ _06562_ _03302_ _03260_ _06565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_158_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10832__I1 mod.u_cpu.rf_ram.memory\[388\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14489_ _00343_ net3 mod.u_cpu.rf_ram.memory\[443\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09159__S _03442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_162_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_255_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14360__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15486__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13917__B _06640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08981_ _01428_ _01429_ _03286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_244_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13534__I0 mod.u_arbiter.i_wb_cpu_dbus_adr\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07932_ _02155_ _02236_ _02239_ _02166_ _02240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_257_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_228_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07863_ _01806_ _02171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_69_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_229_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_244_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09602_ _03757_ _03814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_99_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_216_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07794_ _02057_ _02102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09533_ _03756_ _03757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_243_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08469__A2 _02768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07516__I1 mod.u_cpu.rf_ram.memory\[349\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_184_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_240_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_225_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09464_ _03685_ _03690_ _03691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_227_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__10520__I0 _04469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_227_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__07141__A2 mod.u_cpu.cpu.immdec.imm19_12_20\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08415_ _01459_ _02701_ _02721_ _02722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_09395_ _03631_ _03624_ _03620_ _03632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_178_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_196_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_212_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08346_ _01592_ _02643_ _02652_ _02653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_149_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11599__S _05206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12782__I _05919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_192_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08277_ _01466_ _02038_ _02448_ _02584_ _00000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_20_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12973__B2 _03353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10823__I1 mod.u_cpu.rf_ram.memory\[38\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08641__A2 mod.u_cpu.rf_ram.memory\[172\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14703__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07228_ _01492_ _01536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07159_ _01463_ mod.u_cpu.cpu.immdec.imm19_12_20\[8\] _01467_ mod.u_cpu.cpu.immdec.imm24_20\[4\]
+ _01468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__10587__I0 _04514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_234_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10170_ _01640_ _04229_ _04231_ _00242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_154_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_156_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14853__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07825__B _02132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_247_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_263_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_235_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15209__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13860_ _06465_ _06744_ _06840_ _06854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_41_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12811_ _05630_ _06030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_263_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_216_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13791_ _06791_ _06714_ _06792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_74_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08004__S1 _02295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11861__I _05386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15530_ _01301_ net3 mod.u_cpu.cpu.immdec.imm7 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12742_ _05985_ _01060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_43_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_16_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10511__I0 _04467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07132__A2 _01440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_231_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__14233__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_230_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15359__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15461_ _01235_ net3 mod.u_cpu.cpu.ctrl.o_ibus_adr\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12673_ _05919_ _05940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09409__A1 _03561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11624_ _05222_ mod.u_cpu.rf_ram.memory\[262\]\[0\] _05223_ _05224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__11216__A1 _04668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14412_ _00266_ net3 mod.u_cpu.rf_ram.memory\[481\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12264__I0 _05660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15392_ _01167_ net3 mod.u_cpu.rf_ram.memory\[59\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_129_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11767__A2 _05321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12964__A1 mod.u_cpu.cpu.ctrl.i_iscomp vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09424__A4 _03637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11555_ _05177_ _05178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_14343_ _00197_ net3 mod.u_cpu.rf_ram.memory\[516\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_183_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08391__B _02697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14383__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_155_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10506_ _04442_ _04464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_184_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14274_ _00128_ net3 mod.u_cpu.rf_ram.memory\[550\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_144_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11486_ _03773_ _05132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_13225_ _06331_ _06332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13764__I0 mod.u_cpu.cpu.immdec.imm19_12_20\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10437_ _04272_ _04407_ _04417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_171_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11101__I _04847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12192__A2 _05611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_13156_ _06269_ _01190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_152_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10368_ _04369_ _04335_ _04370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_83_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12107_ _02210_ _05553_ _05554_ _00856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__13229__S _06335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_170_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13087_ _03941_ _06030_ _06227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_239_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10299_ _04322_ _04303_ _04323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_111_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_214_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_12038_ _05508_ _00833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_111_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08699__A2 _03005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_226_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_211_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_266_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_225_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_18_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_13989_ _06942_ _06954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11771__I _03903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_207_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_20_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_222_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_209_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_234_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3090 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10502__I0 _04453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_222_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08320__A1 _02611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_209_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_221_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08200_ mod.u_cpu.rf_ram.memory\[560\]\[0\] mod.u_cpu.rf_ram.memory\[561\]\[0\] mod.u_cpu.rf_ram.memory\[562\]\[0\]
+ mod.u_cpu.rf_ram.memory\[563\]\[0\] _02507_ _02473_ _02508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_33_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_194_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14726__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_178_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09180_ _03461_ _00018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_175_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11758__A2 _05279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_202_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08131_ mod.u_cpu.rf_ram.memory\[47\]\[0\] _02439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_147_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09820__A1 _03870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_179_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08062_ mod.u_cpu.rf_ram.memory\[77\]\[0\] _02370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_107_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14876__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_190_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08387__A1 _02532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13380__A1 _06139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_255_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11946__I _05132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10850__I _04620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_142_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08964_ mod.u_cpu.cpu.mem_bytecnt\[0\] _03269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_103_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08139__A1 _01471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_229_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14180__I0 _07081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07915_ _02066_ mod.u_cpu.rf_ram.memory\[214\]\[0\] _02222_ _01821_ _02223_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_130_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08895_ _02483_ mod.u_cpu.rf_ram.memory\[566\]\[1\] _03201_ _02487_ _03202_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_96_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13683__A2 _06475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_245_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07846_ _01749_ _02154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_83_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14256__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07777_ _02084_ _02085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__11681__I _05262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15501__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09516_ _03739_ _03740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_266_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07114__A2 _01422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08311__A1 _02611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_212_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08195__C _02465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09447_ _03323_ _03324_ _03676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_242_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_213_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_213_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_197_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_240_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09378_ _03610_ _03608_ _03616_ _03617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_197_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_166_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08329_ _02421_ _02635_ _02636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_137_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_193_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11340_ _05032_ mod.u_cpu.rf_ram.memory\[30\]\[1\] _05029_ _05033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_137_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_192_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_158_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_197_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11271_ _04983_ _04984_ _04985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_153_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_238_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08378__A1 _02560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13010_ _06105_ mod.u_cpu.rf_ram.memory\[86\]\[1\] _06175_ _06177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__13371__A1 _06463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10222_ _04268_ _00257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13371__B2 _06466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11856__I _05328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10153_ _04147_ _04217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__15031__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14961_ _00815_ net3 mod.u_cpu.rf_ram.memory\[216\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10084_ _03804_ _04168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_121_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11792__S _05339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13674__A2 _06370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_208_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13912_ _06471_ _06823_ _06390_ _06660_ _06892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__09342__A3 _03586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_208_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14892_ _00746_ net3 mod.u_cpu.rf_ram.memory\[239\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_114_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08550__A1 _01934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_207_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13843_ _06677_ _06838_ _01308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__15181__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_262_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_223_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11437__A1 _04821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14749__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10201__S _04252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13774_ _06289_ _06775_ _06643_ _06317_ _06776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_10986_ _04703_ _04788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_128_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09061__I mod.u_cpu.cpu.csr_imm vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_204_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07736__S0 _02041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_188_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11988__A2 _05475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15513_ _01284_ net3 mod.u_cpu.rf_ram.memory\[329\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_43_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_231_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12725_ _05974_ _01054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_231_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_203_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08853__A2 mod.u_cpu.rf_ram.memory\[38\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_188_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_188_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15444_ _01218_ net3 mod.u_arbiter.i_wb_cpu_ibus_adr\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_157_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12656_ _05918_ mod.u_cpu.rf_ram.memory\[145\]\[0\] _05928_ _05929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_15_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__14899__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_198_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12937__A1 _06057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11607_ _05212_ _00698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_157_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15375_ _01150_ net3 mod.u_cpu.rf_ram.memory\[79\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_141_1243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12587_ _05373_ _05882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_106_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13311__I _06134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14326_ _00180_ net3 mod.u_cpu.rf_ram.memory\[524\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_129_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11538_ _05162_ mod.u_cpu.rf_ram.memory\[277\]\[1\] _05165_ _05167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__11460__I1 mod.u_cpu.rf_ram.memory\[28\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_184_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11469_ _05118_ _05119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_14257_ _00111_ net3 mod.u_cpu.rf_ram.memory\[55\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_7_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08369__A1 _02668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_256_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13208_ _06311_ _06314_ _06315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_125_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07416__I0 mod.u_cpu.rf_ram.memory\[400\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14188_ _03699_ mod.u_cpu.rf_ram.memory\[244\]\[0\] _07089_ _07090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_152_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11766__I _03944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11912__A2 _05423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10670__I _04568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_258_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13139_ mod.u_arbiter.i_wb_cpu_rdt\[21\] mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat\[5\]
+ _06258_ _06260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_98_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10971__I0 _04772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14279__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_239_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_239_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13665__A2 _06659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15524__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08216__S1 _02495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07700_ _01992_ _01996_ _02006_ _02007_ _02008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_227_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08680_ mod.u_cpu.rf_ram.memory\[209\]\[1\] _02987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_39_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_266_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_254_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07631_ mod.u_cpu.rf_ram.memory\[311\]\[0\] _01939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_66_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13417__A2 _04847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07562_ _01550_ _01870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10111__S _04185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_207_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09301_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[12\] _03552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_146_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07493_ mod.u_cpu.rf_ram.memory\[440\]\[0\] mod.u_cpu.rf_ram.memory\[441\]\[0\] mod.u_cpu.rf_ram.memory\[442\]\[0\]
+ mod.u_cpu.rf_ram.memory\[443\]\[0\] _01753_ _01771_ _01801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__08844__A2 _03147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11006__I _04620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09232_ _03492_ _03493_ _03494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_222_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_210_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_222_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_210_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08743__C _02148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12928__A1 _05742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09163_ _03450_ _00012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08114_ mod.u_cpu.rf_ram.memory\[48\]\[0\] mod.u_cpu.rf_ram.memory\[49\]\[0\] mod.u_cpu.rf_ram.memory\[50\]\[0\]
+ mod.u_cpu.rf_ram.memory\[51\]\[0\] _02421_ _02350_ _02422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_119_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_174_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09094_ _03349_ _03395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_162_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_257_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08045_ mod.u_cpu.rf_ram.memory\[69\]\[0\] _02353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_174_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15054__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10167__A1 _03896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_192_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09996_ _03702_ _03939_ _04106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_88_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13105__A1 _04107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08780__A1 _01446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_130_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xtiny_user_project_109 la_data_out[27] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_4505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08947_ _03251_ _03252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_4516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_4527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12703__I1 _05622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_151_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11667__A1 _04226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_151_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08878_ _02592_ _03177_ _03184_ _01836_ _03185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_3826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08532__A1 _02059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_244_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07829_ mod.u_cpu.rf_ram.memory\[167\]\[0\] _02137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_3859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11419__A1 _04539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10840_ _04281_ _04687_ _04688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10021__S _04122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_260_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_198_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10890__A2 _04722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13813__C1 _06812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_198_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_198_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_213_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12092__A1 _05408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_213_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10771_ _04641_ mod.u_cpu.rf_ram.memory\[398\]\[1\] _04638_ _04642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_129_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10956__S _04767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_240_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07194__S1 _01501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12510_ _05827_ mod.u_cpu.rf_ram.memory\[168\]\[0\] _05832_ _05833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_13490_ _03616_ _06551_ _06552_ _03624_ _06553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_139_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08653__C _02139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12441_ _05779_ _00965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_226_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_205_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_201_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08599__A1 _01672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_197_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12372_ _05729_ mod.u_cpu.rf_ram.memory\[499\]\[1\] _05733_ _05735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_15160_ _01013_ net3 mod.u_cpu.rf_ram.memory\[154\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08225__I _02532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_193_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_193_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11787__S _05336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11323_ _05019_ _05020_ _05021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_165_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14111_ _07021_ mod.u_cpu.rf_ram.memory\[87\]\[0\] _07039_ _07040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_180_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15091_ _00945_ net3 mod.u_cpu.rf_ram.memory\[178\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12970__I _03369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_197_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11254_ _04972_ _00585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_14042_ mod.u_arbiter.i_wb_cpu_rdt\[23\] _06987_ _06993_ mod.u_arbiter.i_wb_cpu_dbus_dat\[23\]
+ _06994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_141_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14421__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15547__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10205_ _04249_ mod.u_cpu.rf_ram.memory\[488\]\[0\] _04256_ _04257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_11185_ _04925_ _00563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_133_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10136_ _03866_ _04202_ _04206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_95_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_212_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_209_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_236_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14944_ _00798_ net3 mod.u_cpu.rf_ram.memory\[169\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10067_ _04156_ _00214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__14571__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_208_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_169_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_236_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08523__A1 _01864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_14875_ _00729_ net3 mod.u_cpu.rf_ram.memory\[252\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_263_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13826_ _06471_ _06823_ _06695_ _06490_ _06824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_189_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_91_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10881__A2 _04709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__14072__A2 _07014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13757_ _06492_ _06319_ _06713_ _06744_ _06365_ _06761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_10969_ _04774_ mod.u_cpu.rf_ram.memory\[366\]\[0\] _04776_ _04777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_245_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08382__S0 _02688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12708_ _05962_ _05963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_13688_ _06494_ _06644_ _06696_ _06697_ _06698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_176_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_223_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_15427_ _01202_ net3 mod.u_cpu.rf_ram.memory\[92\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12639_ _05907_ mod.u_cpu.rf_ram.memory\[148\]\[1\] _05915_ _05917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_157_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15077__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_191_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_200_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15358_ _01133_ net3 mod.u_cpu.cpu.genblk3.csr.mcause3_0\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_172_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09251__A2 _03510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10397__A1 _04230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14309_ _00163_ net3 mod.u_cpu.rf_ram.memory\[533\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_171_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15289_ _00048_ net4 mod.u_scanchain_local.module_data_in\[46\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_160_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10149__A1 _01648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_171_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13886__A2 _06285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_252_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09850_ _03945_ _04007_ _04008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_98_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_259_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_213_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__14914__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_213_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08801_ _02204_ mod.u_cpu.rf_ram.memory\[68\]\[1\] _03107_ _03108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_140_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_252_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09781_ _03878_ _03829_ _03955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08732_ mod.u_cpu.rf_ram.memory\[248\]\[1\] mod.u_cpu.rf_ram.memory\[249\]\[1\] mod.u_cpu.rf_ram.memory\[250\]\[1\]
+ mod.u_cpu.rf_ram.memory\[251\]\[1\] _03001_ _01525_ _03039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_6_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08514__A1 _02526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08738__C _01702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08663_ _02711_ _02969_ _02970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_67_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_226_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07614_ _01920_ _01921_ _01922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_208_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08594_ mod.u_cpu.rf_ram.memory\[256\]\[1\] mod.u_cpu.rf_ram.memory\[257\]\[1\] mod.u_cpu.rf_ram.memory\[258\]\[1\]
+ mod.u_cpu.rf_ram.memory\[259\]\[1\] _01837_ _02252_ _02901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_1709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_242_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_183_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08117__I1 _02422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_207_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_263_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07545_ mod.u_cpu.rf_ram.memory\[376\]\[0\] mod.u_cpu.rf_ram.memory\[377\]\[0\] mod.u_cpu.rf_ram.memory\[378\]\[0\]
+ mod.u_cpu.rf_ram.memory\[379\]\[0\] _01837_ _01838_ _01853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__10776__S _04645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08817__A2 _03123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_241_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_222_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11821__A1 _05239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07476_ _01689_ mod.u_cpu.rf_ram.memory\[430\]\[0\] _01781_ _01783_ _01784_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_179_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09490__A2 _03715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_210_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09215_ mod.u_scanchain_local.module_data_in\[34\] mod.u_arbiter.i_wb_cpu_dbus_dat\[29\]
+ _03479_ _03481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_50_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09146_ _03405_ _03439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__12621__I0 _05904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_194_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14444__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09077_ mod.u_cpu.cpu.alu.add_cy_r _03308_ _03379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_190_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_194_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12129__A2 _05568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08028_ _02104_ _02311_ _02335_ _02336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_155_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11188__I0 _04918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10016__S _04119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14594__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5003 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xtiny_user_project_15 io_oeb[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_235_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5014 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_89_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xtiny_user_project_26 io_oeb[18] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_5025 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_162_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_249_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xtiny_user_project_37 io_oeb[29] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__13835__B _06812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5036 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_162_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10560__A1 _04209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtiny_user_project_48 io_out[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_09979_ _04095_ _00187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_5047 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5058 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xtiny_user_project_59 io_out[15] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_5069 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_218_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12990_ _05780_ _06161_ _03373_ _06162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_218_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07308__A2 mod.u_cpu.rf_ram.memory\[510\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_4368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11941_ _05442_ mod.u_cpu.rf_ram.memory\[220\]\[0\] _05444_ _05445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_176_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2900 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10312__A1 _04168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_245_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13126__I _05785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2911 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2922 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14660_ _00514_ net3 mod.u_cpu.rf_ram.memory\[357\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2933 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11872_ _05394_ _00781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2944 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10863__A2 _04704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2955 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_221_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2966 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2977 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13611_ mod.u_cpu.cpu.alu.cmp_r _03687_ _03305_ _06624_ _06630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_26_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10823_ _04663_ mod.u_cpu.rf_ram.memory\[38\]\[0\] _04676_ _04677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08808__A2 _03097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2988 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14591_ _00445_ net3 mod.u_cpu.rf_ram.memory\[392\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2999 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13062__S _06209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13801__A2 _06774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_241_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_201_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13542_ _06583_ _06589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_111_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_242_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10754_ _04630_ _00427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_111_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09481__A2 _01441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_186_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07331__I2 mod.u_cpu.rf_ram.memory\[490\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10485__I _04429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13473_ _06542_ _01234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_10685_ _04315_ _04575_ _04585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_71_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08116__S0 _02242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_200_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15212_ _01065_ net3 mod.u_cpu.rf_ram.memory\[80\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_185_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12424_ _05769_ _00958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_127_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15143_ _00996_ net3 mod.u_cpu.rf_ram.memory\[163\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_154_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12355_ _05713_ mod.u_cpu.rf_ram.memory\[122\]\[0\] _05722_ _05723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07794__I _02057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14937__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13317__A1 _03271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11306_ _05009_ _00600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_12286_ _05662_ mod.u_cpu.rf_ram.memory\[18\]\[0\] _05675_ _05676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_153_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15074_ _00928_ net3 mod.u_cpu.rf_ram.memory\[184\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_153_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11237_ _04960_ _04961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_14025_ mod.u_arbiter.i_wb_cpu_dbus_dat\[20\] _06978_ _06981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_253_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_150_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08744__A1 _02933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11168_ _04913_ _04906_ _04914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_136_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10119_ _04147_ _04193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_110_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11099_ _04867_ _00535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_64_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09514__I _03737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_222_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_14927_ _00781_ net3 mod.u_cpu.rf_ram.memory\[72\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_49_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_209_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_208_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_209_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14317__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14858_ _00712_ net3 mod.u_cpu.rf_ram.memory\[24\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_224_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14045__A2 _06987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13809_ _06401_ _06808_ _06809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_205_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12875__I _06072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14789_ _00643_ net3 mod.u_cpu.rf_ram.memory\[293\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_223_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09847__I1 mod.u_cpu.rf_ram.memory\[542\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_260_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_204_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08355__S0 _02385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07330_ _01637_ _01638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__11803__A1 _04539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_189_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_220_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_220_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_188_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14467__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07261_ _01568_ _01569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_32_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_176_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09000_ mod.u_cpu.cpu.alu.add_cy_r mod.u_cpu.cpu.alu.i_rs1 _03304_ _03305_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_118_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07192_ _01499_ _01500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_157_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07235__A1 _01511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_258_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_145_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_219_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13159__I1 mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08983__A1 mod.u_cpu.cpu.branch_op vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09902_ _04043_ _04044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_193_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_160_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08735__A1 _02179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14108__I0 _07028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_263_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12531__A2 _04528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09833_ _03994_ _03995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_59_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10542__A1 _04352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10393__I1 mod.u_cpu.rf_ram.memory\[460\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_258_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12051__S _05516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09764_ _03941_ _03942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08468__C _01631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08715_ _02027_ _03021_ _03022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_132_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_227_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09695_ _03855_ _03886_ _03887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_132_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08594__S0 _01837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08646_ _01670_ _02945_ _02952_ _02122_ _02953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_70_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10845__A2 _04687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15242__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_187_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_55_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_35 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_70_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_54_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08577_ mod.u_cpu.rf_ram.memory\[280\]\[1\] mod.u_cpu.rf_ram.memory\[281\]\[1\] mod.u_cpu.rf_ram.memory\[282\]\[1\]
+ mod.u_cpu.rf_ram.memory\[283\]\[1\] _02020_ _01995_ _02884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_230_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_161_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13795__B2 _06735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07528_ _01677_ _01836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__12842__I0 _06038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09463__A2 _03276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15392__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07459_ _01751_ _01756_ _01764_ _01766_ _01767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_122_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_210_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10470_ _04439_ _04438_ _04440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_136_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09129_ _03392_ _03426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_159_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12140_ _05387_ _05576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_163_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12770__A2 _05952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10781__A1 _04233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_190_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12071_ _05518_ mod.u_cpu.rf_ram.memory\[63\]\[1\] _05528_ _05530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_46_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08726__A1 _02161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11022_ _04803_ mod.u_cpu.rf_ram.memory\[358\]\[0\] _04813_ _04814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_132_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_133_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08378__C _02594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_206_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12973_ mod.u_cpu.cpu.genblk3.csr.mstatus_mie _06145_ _06148_ _03353_ _06149_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_264_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14712_ _00566_ net3 mod.u_cpu.rf_ram.memory\[331\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_166_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11924_ _05421_ _05432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_206_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_233_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14643_ _00497_ net3 mod.u_cpu.rf_ram.memory\[366\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_233_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11855_ _05382_ _00776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_33_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_205_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07789__I _02096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08394__B _02105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_260_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08337__S0 _02385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10806_ _04665_ _00444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_199_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12833__I0 _06038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14574_ _00428_ net3 mod.u_cpu.rf_ram.memory\[400\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_82_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11786_ _05334_ _05335_ _05336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_13525_ _06577_ _06578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_41_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10737_ _04618_ _00422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_186_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13456_ _06510_ _06531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_10668_ _04560_ mod.u_cpu.rf_ram.memory\[415\]\[1\] _04571_ _04573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_173_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_220_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10943__I _04708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12407_ _05725_ _05757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_177_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_13387_ _06064_ _06482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_10599_ _04514_ mod.u_cpu.rf_ram.memory\[426\]\[1\] _04524_ _04526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_127_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09509__I _03733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10072__I0 _04148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07768__A2 _02075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08965__A1 _03269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15126_ _00979_ net3 mod.u_cpu.rf_ram.memory\[16\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12338_ _05710_ _05711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_181_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_154_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15115__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13010__I0 _06105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15057_ _00911_ net3 mod.u_cpu.rf_ram.memory\[191\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12269_ _05664_ _00908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_142_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08980__A4 _01422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13710__A1 _06694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14008_ _06967_ _06968_ _01343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_123_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10524__A1 _04180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10375__I1 mod.u_cpu.rf_ram.memory\[462\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08812__S1 _02388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09390__A1 _03564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15265__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_233_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_256_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_237_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07940__A2 mod.u_cpu.rf_ram.memory\[236\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_37_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_209_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_209_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13474__B1 _06540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08500_ _02778_ _02799_ _02806_ _01870_ _02807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_09480_ _01461_ _03705_ _03706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_110_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12029__A1 _05239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08431_ _02244_ _02737_ _02738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_252_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_197_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07920__C _01683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07699__I _01787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_205_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13777__A1 _06667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08362_ mod.u_cpu.rf_ram.memory\[485\]\[1\] _02669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_149_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09445__A2 _03674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_177_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07313_ mod.u_cpu.rf_ram.memory\[480\]\[0\] mod.u_cpu.rf_ram.memory\[481\]\[0\] mod.u_cpu.rf_ram.memory\[482\]\[0\]
+ mod.u_cpu.rf_ram.memory\[483\]\[0\] _01605_ _01570_ _01621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_32_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07456__A1 _01689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_220_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08293_ _01607_ _02599_ _02600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_108_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11014__I _04250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_192_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07244_ _01551_ _01552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_30_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_176_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11949__I _05405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_178_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07175_ _01482_ _01483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_192_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10063__I0 _04140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_191_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08708__A1 _02209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_207_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15608__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_143_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08184__A2 _02474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09816_ mod.u_cpu.rf_ram.memory\[545\]\[0\] _03925_ _03981_ _03982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_259_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07931__A2 mod.u_cpu.rf_ram.memory\[230\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_189_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08198__C _02505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09747_ _03733_ _03928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__14632__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_246_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2004 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09133__A1 _03363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2015 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11866__I1 mod.u_cpu.rf_ram.memory\[70\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09678_ _03855_ _03873_ _03874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2026 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_199_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2037 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2048 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08926__C _02539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2059 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_203_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08629_ mod.u_cpu.rf_ram.memory\[180\]\[1\] mod.u_cpu.rf_ram.memory\[181\]\[1\] mod.u_cpu.rf_ram.memory\[182\]\[1\]
+ mod.u_cpu.rf_ram.memory\[183\]\[1\] _02085_ _02086_ _02936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_265_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_215_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_188_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_203_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11125__S _04884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_242_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13768__A1 _03674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11640_ _05234_ mod.u_cpu.rf_ram.memory\[260\]\[1\] _05232_ _05235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__14782__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13768__B2 _06411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07402__I _01509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_243_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07447__A1 _01753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11571_ _05133_ _05188_ _05189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_195_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_211_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13310_ _06403_ _06407_ _06408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_195_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10522_ _04467_ mod.u_cpu.rf_ram.memory\[43\]\[1\] _04473_ _04475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_195_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14290_ _00144_ net3 mod.u_cpu.rf_ram.memory\[542\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_6_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15138__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12464__B _05801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_183_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14193__A1 _07092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13241_ _03771_ _06344_ _06345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10453_ _04251_ _03905_ _04427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_182_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12743__A2 _05552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_123_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10384_ _04230_ _04381_ _04382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_13172_ _06047_ _06279_ _01196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_123_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_163_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12123_ _05559_ mod.u_cpu.rf_ram.memory\[20\]\[0\] _05564_ _05565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_2_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15288__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12054_ _05518_ mod.u_cpu.rf_ram.memory\[61\]\[1\] _05516_ _05519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_151_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_266_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_250_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09372__A1 _03563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11005_ _04801_ _00507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_77_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_238_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_252_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09124__A1 _03392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_265_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11857__I1 mod.u_cpu.rf_ram.memory\[6\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12956_ _06121_ _06130_ _06132_ _06133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__13742__C _06423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_206_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_234_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11907_ _05406_ mod.u_cpu.rf_ram.memory\[224\]\[1\] _05418_ _05420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_3294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12887_ _05896_ _06080_ _06081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_61_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14626_ _00480_ net3 mod.u_cpu.rf_ram.memory\[374\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_60_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11838_ _05370_ _00771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13759__B2 _06475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_199_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_187_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14557_ _00411_ net3 mod.u_cpu.rf_ram.memory\[40\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11769_ mod.u_cpu.rf_ram.memory\[237\]\[1\] _05230_ _05321_ _05324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_159_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13508_ mod.u_cpu.cpu.ctrl.i_jump _03325_ _06563_ _06564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_186_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14488_ _00342_ net3 mod.u_cpu.rf_ram.memory\[443\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10993__A1 _04792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14184__A1 _01985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_179_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13439_ _06521_ _01221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_220_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_179_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13189__C _06285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08938__A1 _01459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14505__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08143__I _02152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_127_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15109_ _00963_ net3 mod.u_cpu.rf_ram.memory\[173\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_170_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08980_ mod.u_cpu.cpu.state.genblk1.misalign_trap_sync_r _03284_ mod.u_cpu.cpu.genblk3.csr.o_new_irq
+ _01422_ _03285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_69_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_170_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07931_ _02179_ mod.u_cpu.rf_ram.memory\[230\]\[0\] _02238_ _02164_ _02239_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_142_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13534__I1 mod.u_arbiter.i_wb_cpu_dbus_adr\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07915__C _01821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14655__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_229_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09363__A1 _03489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07862_ _01741_ _02170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_116_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_217_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09601_ _03813_ _00091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_111_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_257_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_231_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__13933__B _03390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_260_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07793_ _01836_ _02095_ _02100_ _02101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_110_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_228_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13998__A1 mod.u_arbiter.i_wb_cpu_rdt\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09532_ _03753_ _03755_ _03756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_83_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__13998__B2 mod.u_arbiter.i_wb_cpu_dbus_dat\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_266_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09702__I _03807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_266_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09910__I0 _04036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09463_ _03252_ _03276_ _03689_ _03690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_197_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_224_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_184_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08414_ _02609_ _02710_ _02720_ _02721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_197_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09394_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[26\] _03631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_178_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09418__A2 _03615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_240_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07429__A1 _01486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_178_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08345_ _02631_ _02644_ _02651_ _02377_ _02652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__12422__A1 _05312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08276_ _01464_ _01465_ _02522_ _02583_ _02584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_138_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07227_ _01493_ _01502_ _01530_ _01534_ _01535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_180_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07158_ _01449_ _01465_ _01467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__13922__A1 _06166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08053__I _01528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15430__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10587__I1 mod.u_cpu.rf_ram.memory\[428\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_195_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07601__A1 _01874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09729__I0 _03890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15580__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08788__S0 _01636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_232_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_234_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_247_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08937__B _02520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09106__A1 _03398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12810_ _06029_ _01084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_13790_ _06291_ _06791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_170_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09612__I _03821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12459__B _03359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07668__A1 _01739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12741_ _05984_ mod.u_cpu.rf_ram.memory\[209\]\[1\] _05982_ _05985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_216_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07560__C _01867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_256_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_216_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15460_ _01234_ net3 mod.u_cpu.cpu.ctrl.o_ibus_adr\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_163_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12672_ _05939_ _01036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_163_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_204_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_169_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14411_ _00265_ net3 mod.u_cpu.rf_ram.memory\[482\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11623_ _04812_ _05214_ _05223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_179_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15391_ _01166_ net3 mod.u_cpu.rf_ram.memory\[59\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_196_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_169_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10275__I0 _04288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14528__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08093__A1 _02352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12964__A2 _06140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14342_ _00196_ net3 mod.u_cpu.rf_ram.memory\[516\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11554_ _05106_ _05177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_156_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10975__A1 _04377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08391__C _02323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10505_ _04463_ _00345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_239_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_14273_ _00127_ net3 mod.u_cpu.rf_ram.memory\[551\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11485_ _04994_ _05130_ _05131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_156_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13913__A1 _06398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13224_ _06323_ _06326_ _06330_ _06331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_109_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_155_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10436_ _04416_ _00323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_170_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14678__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_170_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09593__A1 _03718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_151_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13155_ mod.u_arbiter.i_wb_cpu_rdt\[28\] mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat\[12\]
+ _06268_ _06269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_3_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10367_ _04066_ _04369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_152_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_88_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12106_ _05488_ _05553_ _05554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_124_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_151_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_257_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10298_ _03796_ _04322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_13086_ _06226_ _01163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_105_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_266_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12037_ mod.u_cpu.rf_ram.memory\[5\]\[1\] _05468_ _05506_ _05508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_78_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_266_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_250_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07307__I _01614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_239_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_253_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_207_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13988_ _06951_ _06953_ _01338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_81_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_230_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_240_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_222_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_207_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12939_ _05781_ _06116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3080 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15303__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_209_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3091 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_234_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_222_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_206_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_248_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13979__I _06910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_222_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14609_ _00463_ net3 mod.u_cpu.rf_ram.memory\[383\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_187_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15589_ _01360_ net3 mod.u_arbiter.i_wb_cpu_dbus_dat\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_261_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_187_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08130_ _02156_ mod.u_cpu.rf_ram.memory\[44\]\[0\] _02437_ _02438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_147_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15453__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09820__A2 _03966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08061_ _01644_ _02369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__14157__A1 _06056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_179_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_134_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13904__A1 _06707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10718__A1 _04180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_192_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_115_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13380__A2 _06475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_170_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_249_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11391__A1 _04784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_216_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08963_ mod.u_cpu.cpu.mem_bytecnt\[1\] _03268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11518__I0 _05144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07645__C _01952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07914_ _02220_ _02221_ _02222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_4709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08894_ _02484_ _03200_ _03201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_57_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07845_ mod.u_cpu.rf_ram.memory\[192\]\[0\] mod.u_cpu.rf_ram.memory\[193\]\[0\] mod.u_cpu.rf_ram.memory\[194\]\[0\]
+ mod.u_cpu.rf_ram.memory\[195\]\[0\] _02151_ _02152_ _02153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__07898__A1 _02202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_217_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_216_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_229_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07776_ _01671_ _02084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_09515_ _03738_ _03739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_140_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_213_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_266_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_213_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_227_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08311__A2 _02614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08048__I _01993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09446_ _03371_ mod.u_cpu.cpu.ctrl.pc_plus_4_cy_r _03675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_197_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_200_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12793__I _06018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09377_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[24\] _03616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_166_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08328_ mod.u_cpu.rf_ram.memory\[501\]\[1\] _02635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_165_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_197_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14820__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_181_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08259_ mod.u_cpu.rf_ram.memory\[535\]\[0\] _02567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__10019__S _04122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_181_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_165_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11270_ _04844_ _04984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__13838__B _03334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_181_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_118_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10221_ _04267_ mod.u_cpu.rf_ram.memory\[486\]\[1\] _04264_ _04268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_165_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14970__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10152_ _04216_ _00239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_106_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_239_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_121_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11509__I0 _05147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14960_ _00814_ net3 mod.u_cpu.rf_ram.memory\[216\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10083_ _04167_ _00219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_94_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13911_ _06641_ _06890_ _06891_ _01323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_87_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_263_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_14891_ _00745_ net3 mod.u_cpu.rf_ram.memory\[238\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_181_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__15326__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_208_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_235_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13842_ mod.u_cpu.cpu.immdec.imm24_20\[0\] _06836_ _06837_ mod.u_cpu.cpu.immdec.imm24_20\[1\]
+ _06838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_114_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_251_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_245_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10488__I _04247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_222_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_13773_ _06309_ _06666_ _06775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10985_ _04787_ _00501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_16_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15512_ _01283_ net3 mod.u_cpu.rf_ram.memory\[329\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_43_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07736__S1 _02043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12724_ mod.u_cpu.rf_ram.memory\[137\]\[1\] _05950_ _05972_ _05974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__14350__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15476__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_204_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15443_ _01217_ net3 mod.u_arbiter.i_wb_cpu_ibus_adr\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_54_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12655_ _05742_ _05920_ _05928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_157_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_169_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11606_ mod.u_cpu.rf_ram.memory\[265\]\[0\] _04954_ _05211_ _05212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08066__A1 _01823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_15374_ _01149_ net3 mod.u_cpu.rf_ram.memory\[107\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_196_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12586_ _05881_ _01008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_184_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14139__A1 _03980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14325_ _00179_ net3 mod.u_cpu.rf_ram.memory\[525\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11537_ _01982_ _05165_ _05166_ _00674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_184_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12208__I _03698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07813__A1 _02110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14256_ _00110_ net3 mod.u_cpu.rf_ram.memory\[55\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_128_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11468_ _03993_ _04701_ _05118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_137_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13207_ _06313_ _06314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08369__A2 _02671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07416__I1 mod.u_cpu.rf_ram.memory\[401\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10419_ _04311_ _04404_ _04405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_14187_ _03842_ _05263_ _07089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_174_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11373__A1 _04369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_174_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11399_ _05071_ mod.u_cpu.rf_ram.memory\[2\]\[0\] _05072_ _05073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_139_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_217_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13138_ _06259_ _01182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_151_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07672__S0 _01957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_217_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_174_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10971__I1 mod.u_cpu.rf_ram.memory\[366\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13069_ _05742_ _06193_ _06215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_78_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12173__I0 _05575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_239_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11920__I0 _05413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07630_ _01825_ _01938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_65_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07561_ _01855_ _01861_ _01868_ _01631_ _01869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_241_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09300_ _03546_ _03550_ _03551_ _00051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_94_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_224_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07492_ _01770_ _01792_ _01799_ _01768_ _01800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_222_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_221_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09231_ _03487_ _03493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_22_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14843__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_179_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_194_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10239__I0 _04267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12928__A2 _04704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09162_ _03449_ mod.u_arbiter.i_wb_cpu_dbus_dat\[7\] _03442_ _03450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_147_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08113_ _01919_ _02421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_163_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_266_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09093_ _03297_ _03394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_163_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14993__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_190_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08044_ _01882_ _02352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_135_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_200_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_163_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07280__A2 _01571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12054__S _05516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13377__C _06472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10167__A2 _04228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08331__I _01537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14223__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15349__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09995_ _04105_ _00193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_5207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_130_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13105__A2 _05640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08780__A2 _03077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08946_ _01421_ _03251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_131_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_218_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_215_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13393__B _06486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_245_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08877_ _02476_ _03180_ _03183_ _02083_ _03184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__11667__A2 _05252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11692__I _05249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_217_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08532__A2 mod.u_cpu.rf_ram.memory\[300\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07828_ _01862_ _02136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__10302__S _04323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14373__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15499__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_204_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07759_ _02042_ _02067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__13813__B1 _06807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08296__A1 _02066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12092__A2 _05543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10770_ _04640_ _04641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_164_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_198_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08934__C _02515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_197_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09429_ _03417_ mod.u_scanchain_local.module_data_in\[68\] _03661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_200_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12440_ _05761_ mod.u_cpu.rf_ram.memory\[172\]\[1\] _05777_ _05779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_139_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13041__A1 _05606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08599__A2 _02905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_201_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12371_ _05734_ _00940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_121_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_219_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14110_ _03823_ _05397_ _07039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11322_ _04995_ _05020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_176_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10650__I0 _04560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_197_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15090_ _00944_ net3 mod.u_cpu.rf_ram.memory\[178\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_176_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14041_ _06970_ _06993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_101_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11253_ _04952_ mod.u_cpu.rf_ram.memory\[322\]\[1\] _04970_ _04972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_4_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10204_ _04255_ _04234_ _04256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10402__I0 _04365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11184_ mod.u_cpu.rf_ram.memory\[333\]\[1\] _04819_ _04923_ _04925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_106_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10135_ _04205_ _00233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_95_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14716__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_209_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14943_ _00797_ net3 mod.u_cpu.rf_ram.memory\[221\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10066_ _04148_ mod.u_cpu.rf_ram.memory\[507\]\[0\] _04155_ _04156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_209_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08523__A2 _02829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14874_ _00728_ net3 mod.u_cpu.rf_ram.memory\[252\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_236_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09072__I _03374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13825_ _06664_ _06823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_169_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_223_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__14866__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11107__I _04024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_189_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10011__I _04050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_250_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13756_ _01479_ _06657_ _06760_ _01299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_91_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__13280__A1 _06377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10968_ _04775_ _04759_ _04776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_62_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_203_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_206_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08844__C _02660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12707_ _05694_ _05962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08382__S1 _02475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_206_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13687_ _06292_ _06485_ _06294_ _06305_ _06697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_189_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11043__S _04828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10899_ _04163_ _04709_ _04729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_15426_ _01201_ net3 mod.u_cpu.rf_ram.memory\[93\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12638_ _05916_ _01025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__14080__I0 _06904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_223_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09787__A1 _03870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15357_ _01132_ net3 mod.u_cpu.cpu.genblk3.csr.mcause3_0\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12569_ _04982_ _05870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_145_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10397__A2 _04390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14308_ _00162_ net3 mod.u_cpu.rf_ram.memory\[533\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_172_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15288_ _00047_ net4 mod.u_scanchain_local.module_data_in\[45\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__14246__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14239_ _00093_ net3 mod.u_cpu.rf_ram.memory\[568\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12394__I0 _05745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08211__A1 _02471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_258_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08800_ _03001_ _03106_ _03107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09780_ _03954_ _00129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__14396__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_230_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07990__I _01744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09183__S _03459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15641__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08731_ _03017_ _03030_ _03037_ _02852_ _03038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_227_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07923__C _01978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_254_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08662_ mod.u_cpu.rf_ram.memory\[223\]\[1\] _02969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_27_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_113_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_215_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07613_ mod.u_cpu.rf_ram.memory\[317\]\[0\] _01921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_96_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08593_ _01979_ _02899_ _01788_ _02900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_81_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_183_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_228_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08117__I2 _02423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07544_ _01851_ _01852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13271__A1 _06367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10085__A1 _04168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_179_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11821__A2 _03829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_179_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07475_ _01782_ _01783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_195_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_195_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13232__I _06338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15021__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09214_ _03480_ _00035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_148_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08326__I _01637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_210_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07230__I _01537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11888__S _05402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09145_ mod.u_arbiter.i_wb_cpu_dbus_dat\[2\] _03438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_108_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08450__A1 _02742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09076_ _03377_ _03378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_190_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15171__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08027_ _01693_ _02322_ _02334_ _02335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_163_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07386__B _01693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14739__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08061__I _01644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5004 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_16 io_oeb[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_5015 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_118_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_27 io_oeb[19] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_5026 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09978_ mod.u_cpu.rf_ram.memory\[521\]\[1\] _03929_ _04093_ _04095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07800__I1 mod.u_cpu.rf_ram.memory\[169\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5037 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12137__I0 _05566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xtiny_user_project_38 io_oeb[30] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_49 io_out[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_5048 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_130_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5059 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08929_ mod.u_cpu.rf_ram.memory\[533\]\[1\] _03236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_4325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12837__A1 _06047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14889__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_183_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10699__I0 _04593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_218_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11940_ _05443_ _05423_ _05444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12311__I _05634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10032__S _04129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_206_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2901 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2912 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13851__B _06844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2923 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11871_ _05383_ mod.u_cpu.rf_ram.memory\[72\]\[1\] _05392_ _05394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_3679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2934 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_205_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2945 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_260_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_169_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2956 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13610_ _03365_ _06625_ _06627_ _06629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__08269__A1 _02551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2967 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10822_ _04511_ _03951_ _04676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_232_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12065__A2 _05525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2978 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_14590_ _00444_ net3 mod.u_cpu.rf_ram.memory\[392\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2989 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09620__I _03827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_214_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08664__C _01703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13541_ _06588_ _01256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_10753_ _04626_ mod.u_cpu.rf_ram.memory\[401\]\[1\] _04628_ _04630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_201_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_158_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10871__I0 _04695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07331__I3 mod.u_cpu.rf_ram.memory\[491\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13472_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[17\] _06538_ _06540_ _03588_ _06542_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_10684_ _04522_ _04584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07492__A2 _01792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14269__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_15211_ _01064_ net3 mod.u_cpu.rf_ram.memory\[199\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08116__S1 _02267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12423_ _05753_ mod.u_cpu.rf_ram.memory\[174\]\[0\] _05768_ _05769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__15514__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11576__A1 _04775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10623__I0 _04537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15142_ _00995_ net3 mod.u_cpu.rf_ram.memory\[163\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12354_ _05452_ _05721_ _05722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_126_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11305_ _05007_ mod.u_cpu.rf_ram.memory\[314\]\[0\] _05008_ _05009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_15073_ _00927_ net3 mod.u_cpu.rf_ram.memory\[179\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12285_ _05563_ _03859_ _05675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_5_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10207__S _04256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14024_ _06979_ _06980_ _01347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_113_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11236_ _04959_ _04960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_136_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10000__A1 _03899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09941__A1 _02552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11167_ _04067_ _04913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_136_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_256_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_171_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10118_ _04192_ _00229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_121_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_212_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_209_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11098_ _04862_ mod.u_cpu.rf_ram.memory\[347\]\[1\] _04865_ _04867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_83_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_49_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_5593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_236_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_76_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14926_ _00780_ net3 mod.u_cpu.rf_ram.memory\[72\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_36_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10049_ _04117_ mod.u_cpu.rf_ram.memory\[510\]\[0\] _04144_ _04145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_4870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_263_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_247_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_14857_ _00711_ net3 mod.u_cpu.rf_ram.memory\[25\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_36_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13253__S _06352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15044__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13808_ _06418_ _06449_ _06807_ _06442_ _06808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_251_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14788_ _00642_ net3 mod.u_cpu.rf_ram.memory\[293\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_50_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12300__I0 _05677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_205_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08574__C _01952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_108_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_204_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13739_ _06713_ _06744_ _06745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_149_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08355__S1 _02633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10676__I _04578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11803__A2 _05279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_232_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_220_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08146__I _02453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07260_ _01497_ _01568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_84_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_220_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__15194__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15409_ _01184_ net3 mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_129_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07191_ _01498_ _01499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11501__S _05140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07985__I _01669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09901_ _03697_ _04043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_160_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_259_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08735__A2 mod.u_cpu.rf_ram.memory\[252\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09832_ _01478_ _03993_ _03994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_140_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08291__S0 _01508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12119__I0 _05550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08749__C _01680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09763_ _03940_ _03941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12819__A1 _03751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13227__I _03502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_227_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08714_ mod.u_cpu.rf_ram.memory\[229\]\[1\] _03021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_255_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08499__A1 _02668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08043__S0 _02349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09694_ _03885_ _03886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_67_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08594__S1 _02252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08645_ _02110_ _02948_ _02951_ _02141_ _02952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_82_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_187_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_242_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_162_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_215_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_214_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_54_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08576_ _01979_ _02875_ _02882_ _01989_ _02883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_26_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_70_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_07527_ _01818_ _01834_ _01835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__09999__A1 _04077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14411__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__15537__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_211_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10853__I0 _04695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_195_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08671__A1 _02606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07458_ _01765_ _01766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_210_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_183_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_22_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_210_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_202_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_194_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07389_ _01633_ _01697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_109_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14561__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09128_ _03416_ _03425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_182_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_191_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_191_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10027__S _04126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09059_ _03315_ _03362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_136_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09816__S _03981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12070_ _05529_ _00844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07609__S0 _01774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13846__B _06840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11021_ _04812_ _04788_ _04813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_104_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_235_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_249_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_238_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07563__C _01870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_213_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_4122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_218_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15067__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12972_ _06142_ _06146_ _06147_ _06145_ _06148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__08034__S0 _01673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_245_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_218_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14711_ _00565_ net3 mod.u_cpu.rf_ram.memory\[332\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11923_ _05431_ _00795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_4199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_261_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14642_ _00496_ net3 mod.u_cpu.rf_ram.memory\[366\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11854_ _05366_ mod.u_cpu.rf_ram.memory\[6\]\[0\] _05381_ _05382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_33_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13235__A1 _03751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_233_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_199_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08337__S1 _02633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10805_ _04663_ mod.u_cpu.rf_ram.memory\[392\]\[0\] _04664_ _04665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_2797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13786__A2 _06774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14573_ _00427_ net3 mod.u_cpu.rf_ram.memory\[401\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_242_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11785_ _05262_ _05335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_159_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13524_ _03923_ _06577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_203_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10736_ _04598_ mod.u_cpu.rf_ram.memory\[403\]\[0\] _04617_ _04618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__14904__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_186_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_13455_ _06530_ _01228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_10667_ _01712_ _04571_ _04572_ _00398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_51_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12406_ _05756_ _00953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_126_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08414__A1 _02609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13386_ _06480_ _06447_ _06481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_126_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10598_ _04525_ _00376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_154_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15125_ _00978_ net3 mod.u_cpu.rf_ram.memory\[459\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_103_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12337_ _05709_ _05710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_138_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11120__I _04620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_15056_ _00910_ net3 mod.u_cpu.rf_ram.memory\[191\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12268_ _05662_ mod.u_cpu.rf_ram.memory\[192\]\[0\] _05663_ _05664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_253_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14007_ _03456_ _06964_ _06958_ mod.u_arbiter.i_wb_cpu_dbus_dat\[14\] _06968_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__09914__A1 _03851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11219_ _04936_ mod.u_cpu.rf_ram.memory\[327\]\[1\] _04946_ _04948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_96_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13710__A2 _06363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12199_ _05616_ _00886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_7_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_209_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_49_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12521__I0 _05827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10288__A1 _04315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14909_ _00763_ net3 mod.u_cpu.rf_ram.memory\[49\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__14434__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12886__I _05396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_224_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_224_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08430_ mod.u_cpu.rf_ram.memory\[407\]\[1\] _02737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_197_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12029__A2 _03851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13226__A1 _06139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_212_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_205_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_260_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08361_ _01960_ _02668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_177_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07312_ _01592_ _01601_ _01619_ _01620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__14584__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_225_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08653__A1 _02135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08292_ mod.u_cpu.rf_ram.memory\[453\]\[1\] _02599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__07456__A2 mod.u_cpu.rf_ram.memory\[422\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_258_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_220_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_149_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_220_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07243_ _01550_ _01551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_137_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10460__A1 _04290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11231__S _04956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_178_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07174_ _01472_ _01473_ _01482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_258_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11260__I0 _04976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11030__I _04531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08708__A2 _03013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11012__I0 _04797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08264__S0 _02450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_232_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12760__I0 _05992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09815_ _03757_ _03980_ _03981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__08479__C _02096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_228_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09746_ _03927_ _00122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08016__S0 _01664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_227_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_223_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12512__I0 _05822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_215_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2005 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09677_ _03872_ _03873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_55_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2016 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_265_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2027 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_215_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2038 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_243_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_160_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10310__S _04328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2049 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08628_ _02090_ _02934_ _02935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_215_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13217__A1 _06321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14927__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_215_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_199_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08559_ _01963_ _02865_ _02866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_243_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11779__A1 _04930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_230_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11570_ _05187_ _05130_ _05188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_74_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08644__A1 _02115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_210_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_168_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10521_ _04474_ _00350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_183_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07839__B _01475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_195_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12464__C _03686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_196_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13240_ _05396_ _06344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_136_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10452_ _04426_ _00329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__14193__A2 _05803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_202_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_100_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_108_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11251__I0 _04961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_182_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_201_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13171_ _03510_ _06278_ _06279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_10383_ _04377_ _04380_ _04381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_124_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14307__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12122_ _05563_ _03843_ _05564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_124_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11875__I _05396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12053_ _05483_ _05518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_111_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_250_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_81_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12751__I0 _05984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11004_ mod.u_cpu.rf_ram.memory\[361\]\[1\] _04661_ _04799_ _04801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_266_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07293__C _01587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14457__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07383__A1 _01688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_266_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_219_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07773__I3 mod.u_cpu.rf_ram.memory\[179\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_206_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12955_ _06131_ _06132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_3240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_206_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_248_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11906_ _05419_ _00790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_209_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13208__A1 _06311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08883__A1 _02456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_179_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12886_ _05396_ _06080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_260_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11837_ _05364_ mod.u_cpu.rf_ram.memory\[228\]\[1\] _05368_ _05370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__13759__A2 _06712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10690__A1 _04457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14625_ _00479_ net3 mod.u_cpu.rf_ram.memory\[375\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_92_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_221_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_199_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_183_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_158_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1893 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08635__A1 _02097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14556_ _00410_ net3 mod.u_cpu.rf_ram.memory\[40\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11768_ _02246_ _05321_ _05323_ _00748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_186_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_202_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10442__A1 _04277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11490__I0 _05128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10954__I _03871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10719_ _04598_ mod.u_cpu.rf_ram.memory\[406\]\[0\] _04606_ _04607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_13507_ mod.u_cpu.cpu.ctrl.i_jump _03296_ _06562_ _06563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_201_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14487_ _00341_ net3 mod.u_cpu.rf_ram.memory\[444\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11699_ _05275_ _00727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_158_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13438_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[4\] _06519_ _06520_ _03520_ _06521_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_228_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_155_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_259_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_155_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13369_ _06464_ _06465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_138_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__15232__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15108_ _00962_ net3 mod.u_cpu.rf_ram.memory\[173\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_114_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11785__I _05262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15039_ _00893_ net3 mod.u_cpu.rf_ram.memory\[198\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_07930_ _01819_ _02237_ _02238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_102_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_111_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07861_ _02150_ _02153_ _02167_ _02168_ _02169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_116_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15382__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_229_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09600_ _03800_ mod.u_cpu.rf_ram.memory\[56\]\[1\] _03811_ _03813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_84_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_256_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07792_ _02097_ _02099_ _02100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_209_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_225_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09531_ _03754_ _03721_ _03755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_37_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07931__C _02164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13998__A2 _06952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_225_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09462_ _03686_ _03687_ _03688_ _03689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_52_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_252_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_08413_ _02539_ _02712_ _02719_ _01678_ _02720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_09393_ _03623_ _03629_ _03630_ _00067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_184_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10808__I0 _04666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08344_ _02597_ _02647_ _02650_ _01651_ _02651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_149_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08626__A1 _01486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12422__A2 _05767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_178_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10433__A1 _04414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_220_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08275_ _01459_ _02558_ _02582_ _02583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_123_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_192_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13240__I _05396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07226_ _01533_ _01534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_138_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_192_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07157_ _01464_ _01465_ _01466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_106_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11933__A1 _05078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_191_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_236_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_266_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13686__A1 _06424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09165__I _03451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12733__I0 _05963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08788__S1 _01638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_259_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_248_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_216_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09729_ _03890_ mod.u_cpu.rf_ram.memory\[555\]\[1\] _03912_ _03914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_210_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12110__A1 _05367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11136__S _04891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12740_ _05937_ _05984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_216_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_203_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10672__A1 _04299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15105__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_242_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12671_ _05938_ mod.u_cpu.rf_ram.memory\[121\]\[1\] _05935_ _05939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_179_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_249_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14410_ _00264_ net3 mod.u_cpu.rf_ram.memory\[482\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11622_ _05221_ _05222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_15390_ _01165_ net3 mod.u_cpu.rf_ram.memory\[103\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_230_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_211_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_196_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10424__A1 _04262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14341_ _00195_ net3 mod.u_cpu.rf_ram.memory\[517\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11553_ _05176_ _00680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_183_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10275__I1 mod.u_cpu.rf_ram.memory\[478\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_211_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_196_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10975__A2 _04780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15255__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10504_ _04450_ mod.u_cpu.rf_ram.memory\[442\]\[1\] _04461_ _04463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_14272_ _00126_ net3 mod.u_cpu.rf_ram.memory\[551\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_13_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11484_ _05119_ _05130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_184_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12177__A1 _05325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13223_ _06329_ _06330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10027__I1 _04111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_183_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13913__A2 _06452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10435_ mod.u_cpu.rf_ram.memory\[453\]\[1\] _04383_ _04413_ _04416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_183_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13154_ _06252_ _06268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__09593__A2 _03806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10366_ _04368_ _00301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_100_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12105_ _03850_ _05552_ _05553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_124_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13085_ _06217_ mod.u_cpu.rf_ram.memory\[104\]\[1\] _06224_ _06226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__13677__A1 _06451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10297_ _04321_ _00279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_78_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09075__I _03334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12036_ _05507_ _00832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09345__A2 _03538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_238_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_226_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_265_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_207_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13987_ mod.u_arbiter.i_wb_cpu_rdt\[9\] _06952_ _06947_ mod.u_arbiter.i_wb_cpu_dbus_dat\[9\]
+ _06953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_207_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13325__I _06421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_262_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3070 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08856__A1 _03151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3081 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12938_ _06115_ _01126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_234_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3092 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_146_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_61_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_261_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12869_ _06035_ mod.u_cpu.rf_ram.memory\[409\]\[0\] _06068_ _06069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_146_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_14608_ _00462_ net3 mod.u_cpu.rf_ram.memory\[383\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_15588_ _01359_ net3 mod.u_arbiter.i_wb_cpu_dbus_dat\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_193_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_187_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10684__I _04522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_174_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14539_ _00393_ net3 mod.u_cpu.rf_ram.memory\[418\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_119_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_187_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08060_ mod.u_cpu.rf_ram.memory\[72\]\[0\] mod.u_cpu.rf_ram.memory\[73\]\[0\] mod.u_cpu.rf_ram.memory\[74\]\[0\]
+ mod.u_cpu.rf_ram.memory\[75\]\[0\] _02366_ _02367_ _02368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__08154__I _02116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14157__A2 mod.u_cpu.cpu.state.o_cnt_r\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12168__A1 _05322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_175_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14622__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12605__S _05893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10718__A2 _04599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_143_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_142_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_255_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_216_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11391__A2 _05058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08962_ mod.u_cpu.cpu.ctrl.pc_plus_offset_cy_r _03266_ _03267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__13668__A1 _06677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14772__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07913_ mod.u_cpu.rf_ram.memory\[215\]\[0\] _02221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_233_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08893_ mod.u_cpu.rf_ram.memory\[567\]\[1\] _03200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_155_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07347__A1 _01591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_190_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07844_ _02126_ _02152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_56_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_257_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07898__A2 _02203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__15128__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07775_ _01785_ _02083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_186_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09514_ _03737_ _03738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_140_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_253_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_224_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09445_ _01451_ _03674_ mod.u_cpu.cpu.o_wen1 vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_13_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_213_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_197_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15278__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_240_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_185_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09376_ _03614_ _03615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_212_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_221_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11454__I0 _05108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08327_ mod.u_cpu.rf_ram.memory\[496\]\[1\] mod.u_cpu.rf_ram.memory\[497\]\[1\] mod.u_cpu.rf_ram.memory\[498\]\[1\]
+ mod.u_cpu.rf_ram.memory\[499\]\[1\] _02632_ _02633_ _02634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__10594__I _04247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_178_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_240_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_193_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_193_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08258_ _02245_ _02566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_153_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12159__A1 _03727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11206__I0 _04938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07209_ _01516_ _01517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_152_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08189_ mod.u_cpu.rf_ram.memory\[573\]\[0\] _02497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_165_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_165_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_35 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10220_ _04266_ _04267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_3_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07836__C _02143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10151_ _04215_ mod.u_cpu.rf_ram.memory\[495\]\[1\] _04213_ _04216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_79_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12314__I _03696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13659__A1 _06371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07408__I _01527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09824__S _03987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10082_ _04157_ mod.u_cpu.rf_ram.memory\[505\]\[1\] _04165_ _04167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_82_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_181_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_43_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_199_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13910_ _03679_ _06649_ _06891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_208_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14890_ _00744_ net3 mod.u_cpu.rf_ram.memory\[238\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_48_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_247_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10893__A1 _04322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13841_ _05787_ _06834_ _06837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__10769__I _04496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13145__I _06252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_210_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_169_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_244_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_13772_ _06773_ _06774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_56_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10984_ _04772_ mod.u_cpu.rf_ram.memory\[364\]\[1\] _04785_ _04787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_216_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13831__A1 _06135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_216_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15511_ _01282_ net3 mod.u_arbiter.i_wb_cpu_dbus_adr\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11693__I0 _05271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12723_ _05973_ _01053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_243_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_231_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12654_ _05927_ _01030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_15442_ _01216_ net3 mod.u_cpu.rf_ram.memory\[339\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_19_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_203_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_169_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11605_ _05078_ _05210_ _05211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_141_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14645__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11445__I0 _05087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_175_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08066__A2 _02373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12585_ _05874_ mod.u_cpu.rf_ram.memory\[157\]\[1\] _05879_ _05881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_15373_ _01148_ net3 mod.u_cpu.rf_ram.memory\[107\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_106_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11536_ _05133_ _05165_ _05166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__14139__A2 _04996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14324_ _00178_ net3 mod.u_cpu.rf_ram.memory\[525\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_102_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_172_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_221_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_176_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13347__B1 _06443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14255_ _00109_ net3 mod.u_cpu.rf_ram.memory\[560\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_139_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11467_ _05117_ _00653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_171_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12425__S _05768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14795__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13206_ _06312_ _06313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_99_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10418_ _03942_ _04335_ _04404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_14186_ _07088_ _01401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_256_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11398_ _04196_ _03975_ _05072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_139_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07577__A1 _01874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12570__A1 _05870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13137_ mod.u_arbiter.i_wb_cpu_rdt\[20\] mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat\[4\]
+ _06258_ _06259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_152_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10349_ _04201_ _04353_ _04357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07672__S1 _01958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_174_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13068_ _06214_ _01157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_215_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12173__I1 mod.u_cpu.rf_ram.memory\[76\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12322__A1 _05037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13256__S _06352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12019_ _05496_ _00826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_152_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_266_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10184__I0 _04215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08621__S0 _02070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09533__I _03756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_253_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07481__C _01788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07560_ _01863_ mod.u_cpu.rf_ram.memory\[382\]\[0\] _01866_ _01867_ _01868_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__08829__A1 _02411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08149__I _01634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15420__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_235_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13822__B2 _06820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_206_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07491_ _01773_ _01795_ _01798_ _01785_ _01799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_61_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07501__A1 _01779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08593__B _01788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09230_ mod.u_arbiter.i_wb_cpu_ibus_adr\[1\] _03492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_94_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_222_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_261_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_203_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09161_ mod.u_arbiter.i_wb_cpu_rdt\[10\] _03449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__15570__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09254__A1 _03506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08112_ mod.u_cpu.rf_ram.memory\[52\]\[0\] mod.u_cpu.rf_ram.memory\[53\]\[0\] mod.u_cpu.rf_ram.memory\[54\]\[0\]
+ mod.u_cpu.rf_ram.memory\[55\]\[0\] _02403_ _02152_ _02420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_33_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09092_ _03362_ _03392_ _03300_ _03279_ _03393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_222_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08043_ mod.u_cpu.rf_ram.memory\[64\]\[0\] mod.u_cpu.rf_ram.memory\[65\]\[0\] mod.u_cpu.rf_ram.memory\[66\]\[0\]
+ mod.u_cpu.rf_ram.memory\[67\]\[0\] _02349_ _02350_ _02351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_134_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09006__A1 _03306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_266_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09708__I _03697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_157_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_170_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09994_ _04091_ mod.u_cpu.rf_ram.memory\[518\]\[1\] _04103_ _04105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_192_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07228__I _01492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08945_ _01440_ _03250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_4507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08876_ _02483_ mod.u_cpu.rf_ram.memory\[558\]\[1\] _03182_ _02487_ _03183_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__13393__C _06487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14518__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08612__S0 _01893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09443__I _03391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08487__C _02453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_229_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07827_ _02134_ _02135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_3839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_151_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14066__A1 mod.u_arbiter.i_wb_cpu_rdt\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_229_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__13113__I0 _06237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_226_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07758_ _01704_ _02066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_72_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14668__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_225_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_213_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07689_ _01960_ _01997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_38_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09428_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[31\] _03657_ _03660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_198_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_241_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_198_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_201_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11427__I0 _05071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09359_ _03489_ _03600_ _03601_ _00061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_100_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13041__A2 _06092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11978__I1 _05468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_240_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12370_ _05731_ mod.u_cpu.rf_ram.memory\[499\]\[0\] _05733_ _05734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_165_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13849__B _06455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_181_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11321_ _03821_ _05019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_197_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10650__I1 mod.u_cpu.rf_ram.memory\[418\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14040_ mod.u_arbiter.i_wb_cpu_dbus_dat\[24\] _06989_ _06992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11252_ _04971_ _00584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_181_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10203_ _03932_ _04255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_175_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10402__I1 mod.u_cpu.rf_ram.memory\[458\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11183_ _04924_ _00562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_238_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07138__I _01446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10134_ _04199_ mod.u_cpu.rf_ram.memory\[498\]\[1\] _04203_ _04205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_122_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13076__S _06219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_251_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_209_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14942_ _00796_ net3 mod.u_cpu.rf_ram.memory\[221\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10065_ _03791_ _04143_ _04155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_48_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15443__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_235_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14873_ _00727_ net3 mod.u_cpu.rf_ram.memory\[254\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_208_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14057__A1 mod.u_arbiter.i_wb_cpu_rdt\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_208_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_251_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_224_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13824_ _06821_ _06822_ _01305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_217_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_169_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_165_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_216_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10618__A1 _04539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_182_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__15593__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13755_ mod.u_cpu.cpu.immdec.imm19_12_20\[8\] _06753_ _06709_ _06759_ _06760_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_10967_ _03884_ _04775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09484__A1 _03707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13280__A2 _03424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_204_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12706_ _05961_ _01048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10094__A2 _04174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_188_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13686_ _06424_ _06682_ _06696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10898_ _04694_ _04728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_148_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15425_ _01200_ net3 mod.u_cpu.rf_ram.memory\[93\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12637_ _05904_ mod.u_cpu.rf_ram.memory\[148\]\[0\] _05915_ _05916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09236__A1 _03414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14080__I1 mod.u_cpu.rf_ram.memory\[299\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15356_ _01131_ net3 mod.u_cpu.cpu.genblk3.csr.mcause31 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_106_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12568_ _05812_ _05869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_157_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11519_ _05154_ _00668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_14307_ _00161_ net3 mod.u_cpu.rf_ram.memory\[534\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_89_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10641__I1 _04396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12499_ _05825_ _00977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_15287_ _00046_ net4 mod.u_scanchain_local.module_data_in\[44\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_156_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09528__I _03751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_236_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_14238_ _00092_ net3 mod.u_cpu.rf_ram.memory\[568\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07476__C _01783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_256_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_217_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14169_ _05780_ _07067_ _07077_ _07078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__08211__A2 _02508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07970__A1 _01791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08730_ _02043_ _03033_ _03036_ _01695_ _03037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_140_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_39_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__12846__A2 _06052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_239_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_187_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_227_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09711__A2 _03897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08661_ _02450_ mod.u_cpu.rf_ram.memory\[220\]\[1\] _02967_ _02968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_39_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14810__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07612_ _01919_ _01920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_208_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08592_ mod.u_cpu.rf_ram.memory\[264\]\[1\] mod.u_cpu.rf_ram.memory\[265\]\[1\] mod.u_cpu.rf_ram.memory\[266\]\[1\]
+ mod.u_cpu.rf_ram.memory\[267\]\[1\] _01802_ _01932_ _02899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_82_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_254_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_241_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_148_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_198_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11657__I0 _05234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07543_ _01850_ _01851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_35_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08117__I3 _02424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_201_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_195_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07474_ _01700_ _01782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_223_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__14960__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_210_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09213_ mod.u_arbiter.i_wb_cpu_rdt\[31\] mod.u_arbiter.i_wb_cpu_dbus_dat\[28\] _03479_
+ _03480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_194_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09227__A1 _03371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11033__I _03959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09144_ _03434_ _03435_ _03437_ _00075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_182_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08770__C _02321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15316__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09075_ _03334_ _03377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_30_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08450__A2 _02756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09438__I _03668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08026_ _02293_ _02324_ _02333_ _02291_ _02334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_190_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_235_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14340__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15466__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5005 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_89_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_17 io_oeb[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_5016 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_130_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xtiny_user_project_28 io_oeb[20] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_104_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09977_ _04094_ _00186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_5027 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xtiny_user_project_39 io_oeb[31] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_5038 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_130_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5049 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_118_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_162_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08928_ mod.u_cpu.rf_ram.memory\[528\]\[1\] mod.u_cpu.rf_ram.memory\[529\]\[1\] mod.u_cpu.rf_ram.memory\[530\]\[1\]
+ mod.u_cpu.rf_ram.memory\[531\]\[1\] _02528_ _02543_ _03235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__10313__S _04332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_264_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_258_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12837__A2 _05788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_217_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08859_ _01471_ _03116_ _03165_ _03166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__14490__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2902 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_233_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2913 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11870_ _05393_ _00780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2924 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2935 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2946 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09901__I _03697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2957 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10821_ _04675_ _00449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_60_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_198_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2968 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13262__A2 mod.u_arbiter.i_wb_cpu_rdt\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2979 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_77_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_214_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13423__I _06509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10752_ _04629_ _00426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_13540_ mod.u_arbiter.i_wb_cpu_dbus_adr\[5\] mod.u_arbiter.i_wb_cpu_dbus_adr\[6\]
+ _06584_ _06588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_197_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_207_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_207_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_200_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_231_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13471_ _06541_ _01233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_71_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_199_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10683_ _04583_ _00403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10871__I1 mod.u_cpu.rf_ram.memory\[382\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15210_ _01063_ net3 mod.u_cpu.rf_ram.memory\[199\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12422_ _05312_ _05767_ _05768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_199_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09769__A2 _03943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08453__S _02125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11576__A2 _05191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15141_ _00994_ net3 mod.u_cpu.rf_ram.memory\[164\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12353_ _05720_ _05721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_166_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13298__C _06395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11304_ _04868_ _04990_ _05008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_15072_ _00926_ net3 mod.u_cpu.rf_ram.memory\[179\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08252__I _02559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12284_ _05674_ _00913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_181_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12525__A1 _05164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14023_ mod.u_arbiter.i_wb_cpu_rdt\[18\] _06976_ _06971_ mod.u_arbiter.i_wb_cpu_dbus_dat\[18\]
+ _06980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_135_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11235_ _03737_ _04959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_141_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14190__S _07089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08824__S0 _02403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12703__S _05959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_214_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10000__A2 _04109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11166_ _04912_ _00557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_110_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14833__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07952__A1 _02175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_212_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10117_ _04178_ mod.u_cpu.rf_ram.memory\[500\]\[1\] _04190_ _04192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_49_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_212_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11097_ _04866_ _00534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_49_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__10139__I0 _04199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09083__I net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14925_ _00779_ net3 mod.u_cpu.rf_ram.memory\[70\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10048_ _03752_ _04143_ _04144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_5594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_248_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_209_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_236_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_224_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13534__S _06584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14856_ _00710_ net3 mod.u_cpu.rf_ram.memory\[25\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_4893 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14983__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_223_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08855__C _02852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13807_ mod.u_arbiter.i_wb_cpu_rdt\[27\] mod.u_arbiter.i_wb_cpu_rdt\[11\] _03509_
+ _06807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_90_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_189_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14787_ _00641_ net3 mod.u_cpu.rf_ram.memory\[294\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11999_ _02221_ _05481_ _05482_ _00820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_44_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_205_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13738_ _06743_ _06744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_147_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_220_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_205_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_220_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_204_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15339__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_177_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13669_ _06658_ _06680_ _06681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_220_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_15408_ _01183_ net3 mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_176_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_192_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07190_ _01497_ _01498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_77_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08590__C _01698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11811__I0 _05342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15339_ _01114_ net3 mod.u_cpu.rf_ram.memory\[96\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_117_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08432__A2 mod.u_cpu.rf_ram.memory\[406\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14363__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15489__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09258__I _03407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13713__B1 _06471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09900_ _03837_ _04033_ _04042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08815__S0 _02366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_258_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08196__A1 _02455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09831_ _03754_ _03992_ _03993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_63_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07943__A1 _02180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08291__S1 _02597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_246_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09762_ _03818_ _03939_ _03940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__12819__A2 _05721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08713_ mod.u_cpu.rf_ram.memory\[224\]\[1\] mod.u_cpu.rf_ram.memory\[225\]\[1\] mod.u_cpu.rf_ram.memory\[226\]\[1\]
+ mod.u_cpu.rf_ram.memory\[227\]\[1\] _01507_ _01763_ _03020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_09693_ _03884_ _03885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13952__B _03438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08043__S1 _02350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_265_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08644_ _02115_ mod.u_cpu.rf_ram.memory\[174\]\[1\] _02950_ _01771_ _02951_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_2209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_227_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_55_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10550__I0 _04481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_54_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_199_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_82_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08575_ _01981_ _02878_ _02881_ _01972_ _02882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_1519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__09448__A1 _03334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_35_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_81_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_165_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07526_ _01822_ _01824_ _01829_ _01831_ _01832_ _01833_ _01834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_223_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09999__A2 _04108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_211_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10302__I0 _04313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08120__A1 _02406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11899__S _05414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_211_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07457_ _01527_ _01765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_211_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_211_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14706__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07388_ _01695_ _01696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_176_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09127_ mod.u_arbiter.i_wb_cpu_rdt\[1\] _03424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_176_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_194_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08072__I _01485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09058_ _03306_ _03360_ _03346_ _03361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_159_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_191_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14856__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08009_ mod.u_cpu.rf_ram.memory\[127\]\[0\] _02317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_123_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07609__S1 _01916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13180__A1 _05783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11020_ _03949_ _04812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_173_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_238_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_106_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_265_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_213_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11869__I0 _05385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_181_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_3411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12971_ mod.u_cpu.cpu.genblk3.csr.mstatus_mpie _06142_ _06147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_85_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08034__S1 _01666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14710_ _00564_ net3 mod.u_cpu.rf_ram.memory\[332\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11922_ _05426_ mod.u_cpu.rf_ram.memory\[222\]\[1\] _05429_ _05431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_3444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_206_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_205_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09631__I _03836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_260_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__14236__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14641_ _00495_ net3 mod.u_cpu.rf_ram.memory\[367\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11853_ _05239_ _03951_ _05381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_3499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13235__A2 _06193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10804_ _04255_ _04648_ _04664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08247__I _02308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14572_ _00426_ net3 mod.u_cpu.rf_ram.memory\[401\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11784_ _03917_ _05334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_2798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08111__A1 _01693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07151__I _01439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_214_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07545__S0 _01837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_202_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_201_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13523_ _06576_ _01250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_10735_ _04352_ _04599_ _04617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11602__S _05206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14386__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_220_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15631__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_13454_ _03547_ _06525_ _06526_ _03552_ _06530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_10666_ _04542_ _04571_ _04572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_174_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12405_ _05745_ mod.u_cpu.rf_ram.memory\[176\]\[1\] _05754_ _05756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_13385_ _06397_ _06129_ _06480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_173_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09611__A1 _03818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10597_ _04523_ mod.u_cpu.rf_ram.memory\[426\]\[0\] _04524_ _04525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_127_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_15124_ _00977_ net3 mod.u_cpu.rf_ram.memory\[459\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12336_ _05105_ _05709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_115_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12267_ _05417_ _05650_ _05663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_15055_ _00909_ net3 mod.u_cpu.rf_ram.memory\[192\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_107_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_218_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13171__A1 _03510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11218_ _04947_ _00574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_14006_ mod.u_arbiter.i_wb_cpu_dbus_dat\[15\] _06966_ _06967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09914__A2 _04038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12198_ mod.u_cpu.rf_ram.memory\[201\]\[0\] _05437_ _05615_ _05616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07754__C _01818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_256_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_150_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11149_ _04882_ _04901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_1_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_228_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15011__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_163_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07326__I _01633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_255_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_209_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_5380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_252_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11485__A1 _04994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14908_ _00762_ net3 mod.u_cpu.rf_ram.memory\[49\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_64_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_209_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08585__C _02007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14839_ _00693_ net3 mod.u_cpu.rf_ram.memory\[268\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__15161__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_212_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13226__A2 _06332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_251_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08360_ mod.u_cpu.rf_ram.memory\[480\]\[1\] mod.u_cpu.rf_ram.memory\[481\]\[1\] mod.u_cpu.rf_ram.memory\[482\]\[1\]
+ mod.u_cpu.rf_ram.memory\[483\]\[1\] _01963_ _02666_ _02667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__14729__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08157__I _01747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07311_ _01602_ _01606_ _01617_ _01618_ _01619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_60_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12985__A1 _06113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08291_ mod.u_cpu.rf_ram.memory\[448\]\[1\] mod.u_cpu.rf_ram.memory\[449\]\[1\] mod.u_cpu.rf_ram.memory\[450\]\[1\]
+ mod.u_cpu.rf_ram.memory\[451\]\[1\] _01508_ _02597_ _02598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_149_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09850__A1 _03945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07242_ mod.u_cpu.raddr\[3\] _01550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_177_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12737__A1 _03865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14879__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_1281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_118_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_192_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07173_ _01478_ _01479_ _01480_ _01481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__12407__I _05725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10599__I0 _04514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_259_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09716__I _03903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_236_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07916__A1 _01651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08264__S1 _02451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09814_ _03979_ _03980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_98_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_247_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10771__I0 _04641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14259__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09745_ mod.u_cpu.rf_ram.memory\[553\]\[0\] _03925_ _03926_ _03927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10798__S _04659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08016__S1 _02323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11981__I _05422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15504__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_228_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2006 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09676_ _03871_ _03872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2017 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2028 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_242_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2039 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_215_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08627_ mod.u_cpu.rf_ram.memory\[176\]\[1\] mod.u_cpu.rf_ram.memory\[177\]\[1\] mod.u_cpu.rf_ram.memory\[178\]\[1\]
+ mod.u_cpu.rf_ram.memory\[179\]\[1\] _02048_ _02086_ _02934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_1316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08892__A2 mod.u_cpu.rf_ram.memory\[564\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12276__I0 _05662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_230_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08558_ mod.u_cpu.rf_ram.memory\[309\]\[1\] _02865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_74_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07509_ _01656_ _01816_ _01817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_167_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08489_ _02778_ _02788_ _02795_ _02677_ _02796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__12518__S _05835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_51_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_167_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07298__I3 mod.u_cpu.rf_ram.memory\[507\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10520_ _04469_ mod.u_cpu.rf_ram.memory\[43\]\[0\] _04473_ _04474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_161_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_202_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_202_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10451_ _04410_ mod.u_cpu.rf_ram.memory\[450\]\[1\] _04424_ _04426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_182_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13170_ _03492_ _03412_ _03400_ _06278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_10382_ _04225_ _04379_ _04380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_184_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12121_ _04982_ _05563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_163_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_237_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_191_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__15034__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12052_ _05517_ _00838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_137_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_266_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_238_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11003_ _04800_ _00506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_46_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_266_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_266_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08580__A1 _01998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07383__A2 _01690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_237_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15184__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12954_ _06125_ _06128_ _06131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_3241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_261_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11905_ _05413_ mod.u_cpu.rf_ram.memory\[224\]\[0\] _05418_ _05419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_3274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_234_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13208__A2 _06314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12885_ _06079_ _01109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_233_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_206_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14624_ _00478_ net3 mod.u_cpu.rf_ram.memory\[375\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11836_ _05369_ _00770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10690__A2 _04575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_183_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12967__A1 _03338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14555_ _00409_ net3 mod.u_cpu.rf_ram.memory\[410\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11767_ _05322_ _05321_ _05323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09832__A1 _01478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1894 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_187_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_147_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13506_ _06142_ _03250_ _06562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10718_ _04180_ _04599_ _04606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_14486_ _00340_ net3 mod.u_cpu.rf_ram.memory\[444\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11698_ _05271_ mod.u_cpu.rf_ram.memory\[254\]\[1\] _05273_ _05275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_158_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13437_ _06513_ _06520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_10649_ _04497_ _04560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13392__A1 _06470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_259_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13368_ _06388_ _06464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_155_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15107_ _00961_ net3 mod.u_cpu.rf_ram.memory\[439\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12163__S _05590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12319_ _05698_ _00924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_181_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13299_ _06328_ _06397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09199__I0 mod.u_arbiter.i_wb_cpu_rdt\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_244_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_15038_ _00892_ net3 mod.u_cpu.rf_ram.memory\[198\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_170_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14401__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15527__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_257_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07860_ _01586_ _02168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_69_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_229_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10753__I0 _04626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_3_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07791_ mod.u_cpu.rf_ram.memory\[188\]\[0\] mod.u_cpu.rf_ram.memory\[189\]\[0\] mod.u_cpu.rf_ram.memory\[190\]\[0\]
+ mod.u_cpu.rf_ram.memory\[191\]\[0\] _02092_ _02098_ _02099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_49_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09530_ _03716_ _03717_ _03754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__14551__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08323__A1 _02039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_224_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_188_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09461_ _03681_ _03679_ _03688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_37_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_225_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08412_ _02654_ _02715_ _02718_ _01992_ _02719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_197_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09392_ _03496_ mod.u_scanchain_local.module_data_in\[62\] _03630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_52_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_178_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08343_ _02638_ mod.u_cpu.rf_ram.memory\[510\]\[1\] _02649_ _01821_ _02650_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__09823__A1 _03767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_225_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11630__A1 _04817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08274_ _02571_ _02581_ _02520_ _02582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__10433__A2 _04413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_203_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13758__I0 mod.u_arbiter.i_wb_cpu_rdt\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13907__B1 _06682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07225_ _01532_ _01533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_20_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11041__I _04802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15057__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13383__A1 _03665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_180_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07156_ _01438_ _01465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11233__I1 _04819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12430__I0 _05761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11933__A2 _05438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07988__I1 mod.u_cpu.rf_ram.memory\[105\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13686__A2 _06682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_232_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_219_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07989_ _02091_ _02297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_235_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_228_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09728_ _03913_ _00118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_132_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10321__S _04336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_210_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_216_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12110__A2 _05543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_243_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_167_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09659_ _03858_ _03859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_215_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_216_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_203_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10672__A2 _04575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12670_ _05937_ _05938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_243_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11621_ _04959_ _05221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14340_ _00194_ net3 mod.u_cpu.rf_ram.memory\[517\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11552_ _05159_ mod.u_cpu.rf_ram.memory\[274\]\[0\] _05175_ _05176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_196_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09290__A2 _03538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10503_ _04462_ _00344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_11483_ _05129_ _00657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_14271_ _00125_ net3 mod.u_cpu.rf_ram.memory\[552\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_156_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12177__A2 _05568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13222_ _06328_ _06129_ _06329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_10434_ _01512_ _04413_ _04415_ _00322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_109_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14424__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__13079__S _06219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13153_ _06267_ _01189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_151_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_124_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10365_ _04363_ mod.u_cpu.rf_ram.memory\[464\]\[1\] _04366_ _04368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_87_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12104_ _05432_ _05552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_135_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13084_ _06225_ _01162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_10296_ _04313_ mod.u_cpu.rf_ram.memory\[475\]\[1\] _04319_ _04321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_250_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_239_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_12035_ mod.u_cpu.rf_ram.memory\[5\]\[0\] _05437_ _05506_ _05507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_2_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12724__I1 _05950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_266_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14574__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_215_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08553__A1 _01949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_77_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_266_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_226_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11327__S _05021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_266_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13986_ _06937_ _06952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_93_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09091__I mod.u_cpu.cpu.bufreg.lsb\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_248_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_206_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3060 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12937_ _06057_ _06114_ _06115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_3071 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11160__I0 _04896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_234_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__15821__I net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3082 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3093 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_185_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12868_ _05896_ _04687_ _06068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_222_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_178_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14607_ _00461_ net3 mod.u_cpu.rf_ram.memory\[384\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_221_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11819_ _05350_ mod.u_cpu.rf_ram.memory\[230\]\[1\] _05356_ _05358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_187_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15587_ _01358_ net3 mod.u_arbiter.i_wb_cpu_dbus_dat\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_15_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12799_ _06019_ mod.u_cpu.rf_ram.memory\[12\]\[1\] _06021_ _06023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_1691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_222_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_187_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_159_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14538_ _00392_ net3 mod.u_cpu.rf_ram.memory\[418\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_109_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_230_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_175_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07292__A1 _01505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14469_ _00323_ net3 mod.u_cpu.rf_ram.memory\[453\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_175_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12168__A2 _05595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_190_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_161_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_143_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14917__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_192_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_170_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08170__I _02477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_170_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08961_ mod.u_arbiter.i_wb_cpu_ibus_adr\[0\] _03265_ _03266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_170_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07912_ _01519_ _02220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_233_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08892_ _02478_ mod.u_cpu.rf_ram.memory\[564\]\[1\] _03198_ _03199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_151_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08544__A1 _02295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07843_ _01856_ _02151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_84_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_256_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07774_ _02080_ _02081_ _02082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09513_ _03695_ _03737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_25_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_225_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11151__I0 _04901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_266_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_252_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09444_ _03353_ _03673_ _03674_ mod.u_cpu.cpu.o_wen0 vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_262_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_213_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_80_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09375_ _03486_ _03614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13251__I _06204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_240_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_166_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08326_ _01637_ _02633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_166_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12651__I0 _05918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14447__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_177_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08257_ _02527_ mod.u_cpu.rf_ram.memory\[532\]\[0\] _02564_ _02565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_21_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_229_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12159__A2 _04379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07208_ _01515_ _01516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_119_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08188_ mod.u_cpu.rf_ram.memory\[568\]\[0\] mod.u_cpu.rf_ram.memory\[569\]\[0\] mod.u_cpu.rf_ram.memory\[570\]\[0\]
+ mod.u_cpu.rf_ram.memory\[571\]\[0\] _02494_ _02495_ _02496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_193_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12403__I0 _05753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07139_ _01439_ _01448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_106_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_238_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09176__I _03451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14597__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08783__A1 _02051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08080__I _02126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10150_ _04177_ _04215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_161_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10081_ _04166_ _00218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_173_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_248_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09583__I0 _03740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11147__S _04898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13426__I _06512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13840_ _06835_ _06836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10893__A2 _04709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07424__I _01614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_216_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_249_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_261_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_13771_ _06415_ _06772_ _06773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__11142__I0 _04896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10983_ _04786_ _00500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_167_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15510_ _01281_ net3 mod.u_arbiter.i_wb_cpu_dbus_adr\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_231_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12722_ mod.u_cpu.rf_ram.memory\[137\]\[0\] _05971_ _05972_ _05973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__15222__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12890__I0 _06070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08683__C _02591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15441_ _01215_ net3 mod.u_cpu.rf_ram.memory\[339\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_203_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_128_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12653_ _05923_ mod.u_cpu.rf_ram.memory\[146\]\[1\] _05925_ _05927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_90_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_180_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_230_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11604_ _03723_ _04779_ _05210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_168_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15372_ _01147_ net3 mod.u_cpu.rf_ram.memory\[83\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12584_ _05880_ _01007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_129_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14323_ _00177_ net3 mod.u_cpu.rf_ram.memory\[526\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_23_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15372__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11535_ _05164_ _05130_ _05165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_184_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13347__A1 _06442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13347__B2 _06382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14254_ _00108_ net3 mod.u_cpu.rf_ram.memory\[560\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_172_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11466_ _05108_ mod.u_cpu.rf_ram.memory\[288\]\[1\] _05115_ _05117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_183_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13898__A2 _06881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13205_ mod.u_arbiter.i_wb_cpu_rdt\[8\] mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat\[8\]
+ _03499_ _06312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_143_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10417_ _04403_ _00317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_14185_ _07081_ mod.u_cpu.rf_ram.memory\[279\]\[1\] _07086_ _07088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_11397_ _05045_ _05071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_178_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_125_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10226__S _04269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_180_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10956__I0 _04753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09086__I _03386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08774__A1 _02477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14147__I0 _07055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13136_ _06252_ _06258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__12570__A2 _04913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10348_ _04356_ _00295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10279_ _04308_ _04309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_13067_ _06199_ mod.u_cpu.rf_ram.memory\[106\]\[1\] _06212_ _06214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_140_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_239_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08526__A1 _01872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12018_ _05470_ mod.u_cpu.rf_ram.memory\[214\]\[0\] _05495_ _05496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_79_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_238_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08621__S1 _02071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_266_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_254_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_171_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_207_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13780__B _06380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12086__A1 _04973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08829__A2 _03135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13969_ _06936_ _06939_ _01333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_81_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13822__A2 _06815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_253_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_234_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07490_ _01689_ mod.u_cpu.rf_ram.memory\[438\]\[0\] _01797_ _01763_ _01798_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_263_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_263_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_250_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07501__A2 _01808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15639_ _01410_ net3 mod.u_cpu.cpu.mem_bytecnt\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_34_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_181_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_226_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09160_ _03448_ _00011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_222_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08165__I _02388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_187_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08111_ _01693_ _02392_ _02418_ _02380_ _02419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_148_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09091_ mod.u_cpu.cpu.bufreg.lsb\[1\] _03392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_266_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_175_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11520__S _05153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_175_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09197__S _03469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08042_ _01637_ _02350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_175_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13889__A2 _06836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_200_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10947__I0 _04756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_192_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08765__A1 _02297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10572__A1 _04218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09993_ _04104_ _00192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_142_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_5209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08944_ _03249_ _00002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09724__I _03909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08768__C _02306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_130_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08875_ _02484_ _03181_ _03182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_56_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_257_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08612__S1 _02054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12150__I _05549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07826_ _01634_ _02134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_85_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15245__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07244__I _01551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07757_ _01849_ _02064_ _02065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_198_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_253_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12872__I0 _06070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07688_ mod.u_cpu.rf_ram.memory\[280\]\[0\] mod.u_cpu.rf_ram.memory\[281\]\[0\] mod.u_cpu.rf_ram.memory\[282\]\[0\]
+ mod.u_cpu.rf_ram.memory\[283\]\[0\] _01994_ _01995_ _01996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_129_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15395__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09427_ mod.u_arbiter.i_wb_cpu_dbus_adr\[31\] _03659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_240_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_212_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_197_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12624__I0 _05907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09358_ _03554_ mod.u_scanchain_local.module_data_in\[57\] _03555_ mod.u_arbiter.i_wb_cpu_dbus_adr\[20\]
+ _03601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_166_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07256__A1 _01545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08309_ _02532_ _02615_ _02616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_100_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09289_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[9\] _03542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_166_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13329__A1 _06425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11320_ _05018_ _00605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_153_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_154_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_197_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11251_ _04961_ mod.u_cpu.rf_ram.memory\[322\]\[0\] _04970_ _04971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_107_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10202_ _04254_ _00251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_11182_ mod.u_cpu.rf_ram.memory\[333\]\[0\] _04658_ _04923_ _04924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_136_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_134_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_192_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_171_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10133_ _04204_ _00232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_122_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08508__A1 _02668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09556__I0 _03764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08678__C _01632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14941_ _00795_ net3 mod.u_cpu.rf_ram.memory\[222\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10064_ _04154_ _00213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11363__I0 _05046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_236_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_236_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14872_ _00726_ net3 mod.u_cpu.rf_ram.memory\[254\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_75_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_236_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_76_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07154__I _01462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14057__A2 _06998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12068__A1 _04294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13823_ mod.u_cpu.cpu.immdec.imm30_25\[3\] _06773_ _06812_ mod.u_cpu.cpu.immdec.imm30_25\[4\]
+ _06822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_91_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_217_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12995__I _03686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14188__S _07089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14612__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_235_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13804__A2 _06714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_216_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_204_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_216_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13754_ _06432_ _06755_ _06758_ _06065_ _06759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__10618__A2 _04447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10966_ _04694_ _04774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_232_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_206_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12705_ mod.u_cpu.rf_ram.memory\[13\]\[1\] _05950_ _05959_ _05961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_245_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13685_ _06694_ _06398_ _06695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_70_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10897_ _04727_ _00473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_15424_ _01199_ net3 mod.u_cpu.rf_ram.memory\[94\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_231_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14762__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_188_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12636_ _05535_ _05900_ _05915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_169_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_223_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_15355_ _01130_ net3 mod.u_cpu.cpu.genblk3.csr.mstatus_mpie vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12567_ _05868_ _01002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13759__C _06412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_200_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_200_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14306_ _00160_ net3 mod.u_cpu.rf_ram.memory\[534\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11518_ _05144_ mod.u_cpu.rf_ram.memory\[280\]\[0\] _05153_ _05154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_172_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15286_ _00045_ net4 mod.u_scanchain_local.module_data_in\[43\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_144_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12498_ _05813_ mod.u_cpu.rf_ram.memory\[459\]\[0\] _05824_ _05825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__15118__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12918__I1 _06005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14237_ _00091_ net3 mod.u_cpu.rf_ram.memory\[56\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_109_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11449_ _05104_ _00648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_172_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08747__A1 _02156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07329__I _01568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13740__A1 _06470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09745__S _03926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14168_ _05790_ _06166_ _03393_ _07073_ _07077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_112_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13119_ _06247_ _01175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15268__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14099_ _07032_ _01370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09544__I _03756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_252_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07492__C _01768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_239_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10306__A1 _04163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_230_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_152_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08660_ _02656_ _02966_ _02967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_94_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_215_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__14292__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07611_ _01743_ _01919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_26_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08591_ _02759_ _02894_ _02897_ _02764_ _02898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__14098__S _07030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11515__S _05150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_223_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07542_ _01490_ _01850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11657__I1 mod.u_cpu.rf_ram.memory\[258\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_207_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09475__A2 _03700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07473_ _01779_ _01780_ _01781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07486__A1 _01774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_223_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_222_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09212_ _03414_ _03479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__09227__A2 _03489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09143_ mod.u_arbiter.i_wb_cpu_rdt\[4\] _03436_ _03437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_33_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08986__A1 _03289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_175_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_147_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09074_ _03370_ _03376_ mod.u_cpu.cpu.o_wdata1 vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_148_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_194_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_159_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08025_ _02325_ _02328_ _02332_ _01717_ _02333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_200_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_159_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13031__I0 _06186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_190_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_190_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08738__A1 _02632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13731__A1 mod.u_cpu.cpu.immdec.imm19_12_20\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08779__B _03085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07410__A1 _01703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5006 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_104_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09976_ mod.u_cpu.rf_ram.memory\[521\]\[0\] _03925_ _04093_ _04094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_5017 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xtiny_user_project_18 io_oeb[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_162_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5028 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xtiny_user_project_29 io_oeb[21] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_83_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5039 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08498__C _02453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08927_ _02523_ _03226_ _03233_ _02505_ _03234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_4305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_190_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11345__I0 _05032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14635__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_218_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_4327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_218_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08858_ _01475_ _03141_ _03164_ _03165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_3626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2903 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07809_ mod.u_cpu.rf_ram.memory\[175\]\[0\] _02117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_211_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2914 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2925 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08789_ _01493_ _03095_ _01534_ _03096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_217_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2936 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13798__A1 _06401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2947 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10820_ _04666_ mod.u_cpu.rf_ram.memory\[390\]\[1\] _04673_ _04675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_198_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14785__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2958 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2969 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_77_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07702__I _01581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_198_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10751_ _04622_ mod.u_cpu.rf_ram.memory\[401\]\[0\] _04628_ _04629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_111_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_241_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11224__I _04795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_198_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_213_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13470_ _03578_ _06538_ _06540_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[17\] _06541_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_51_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10682_ _04579_ mod.u_cpu.rf_ram.memory\[413\]\[1\] _04581_ _04583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_199_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12421_ _05725_ _05767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12222__A1 _05019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_224_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_200_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_166_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15140_ _00993_ net3 mod.u_cpu.rf_ram.memory\[164\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_138_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12352_ _05629_ _05720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_127_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13970__A1 _03412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_181_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11303_ _04960_ _05007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13022__I0 _06184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15071_ _00925_ net3 mod.u_cpu.rf_ram.memory\[189\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_153_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12283_ _05660_ mod.u_cpu.rf_ram.memory\[190\]\[1\] _05672_ _05674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_153_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08729__A1 _02632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07149__I _01457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13722__A1 _06463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15410__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14022_ mod.u_arbiter.i_wb_cpu_dbus_dat\[19\] _06978_ _06979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09777__I0 _03916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12525__A2 _04302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11234_ _04958_ _00579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_106_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08824__S1 _02367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08689__B _02995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10387__I1 _04383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11165_ _04896_ mod.u_cpu.rf_ram.memory\[336\]\[1\] _04910_ _04912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_96_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10116_ _04191_ _00228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_251_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11096_ _04864_ mod.u_cpu.rf_ram.memory\[347\]\[0\] _04865_ _04866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_5540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_209_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11336__I0 _05028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_5551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_5562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15560__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14924_ _00778_ net3 mod.u_cpu.rf_ram.memory\[70\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10047_ _04142_ _04143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_5584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_4883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14855_ _00709_ net3 mod.u_cpu.rf_ram.memory\[260\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_5_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_264_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4894 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_236_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_224_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_217_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_205_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13806_ _06735_ _06802_ _06805_ _06332_ _06806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_90_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14786_ _00640_ net3 mod.u_cpu.rf_ram.memory\[294\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_56_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11998_ _05448_ _05481_ _05482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__07612__I _01919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07468__A1 _01774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_232_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13737_ _06288_ _06667_ _06669_ _06743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_72_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_204_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12461__A1 _03359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10949_ _04511_ _03961_ _04763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_189_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13668_ _06677_ _06679_ _06680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_143_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__14202__A2 _06151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15407_ _01182_ net3 mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_12619_ _05886_ _05904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07768__B _01602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13599_ _03694_ _06573_ _06620_ _03659_ _01282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_118_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14508__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09539__I _03761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13961__A1 mod.u_arbiter.i_wb_cpu_rdt\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15338_ _01113_ net3 mod.u_cpu.rf_ram.memory\[98\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11811__I1 mod.u_cpu.rf_ram.memory\[49\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10775__A1 _04643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_219_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07640__A1 _01643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_15269_ _00026_ net4 mod.u_arbiter.i_wb_cpu_rdt\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__13013__I0 _06107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15090__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13713__A1 mod.u_cpu.cpu.immdec.imm19_12_20\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12516__A2 _05835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13713__B2 _06693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08815__S1 _02367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14658__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08196__A2 _02499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09830_ _03806_ _03992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_28_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09761_ _03746_ _03938_ _03939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_258_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11327__I0 _05014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11309__I _04989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08111__C _02380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08712_ _03017_ _03018_ _01870_ _03019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09692_ _03856_ _03883_ _03884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_230_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_227_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_187_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08643_ _02116_ _02949_ _02950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_94_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_215_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11245__S _04966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_254_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_70_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08574_ _01697_ mod.u_cpu.rf_ram.memory\[278\]\[1\] _02880_ _01952_ _02881_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_148_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__09448__A2 _03668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07522__I _01820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_63_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07525_ _01679_ _01833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_39_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07459__A1 _01751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_223_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_228_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_194_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07456_ _01689_ mod.u_cpu.rf_ram.memory\[422\]\[0\] _01761_ _01763_ _01764_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_210_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_241_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07387_ _01491_ _01695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_157_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10066__I0 _04148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_182_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15433__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09126_ _03423_ _00041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__08353__I _01679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10766__A1 _04218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_194_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_191_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09057_ _03355_ mod.u_cpu.cpu.csr_imm _03358_ _03359_ _03360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_68_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12804__S _06024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_237_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13704__A1 _06470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08008_ _01924_ _02316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_190_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__15583__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13180__A2 mod.u_arbiter.i_wb_cpu_rdt\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09959_ _04082_ _00180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_77_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_264_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12970_ _03369_ _06146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_4146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13862__C _06704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09912__I _03738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07698__A1 _01997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11921_ _05430_ _00794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_206_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12691__A1 _03723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14640_ _00494_ net3 mod.u_cpu.rf_ram.memory\[367\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_61_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11852_ _05380_ _00775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_233_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_221_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_199_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10803_ _04621_ _04663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_199_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14571_ _00425_ net3 mod.u_cpu.rf_ram.memory\[402\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_82_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11783_ _05333_ _00753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08972__B _03276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_207_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08111__A2 _02392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_199_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13522_ _03426_ _06575_ _06570_ _06576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07545__S1 _01838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10734_ _04616_ _00421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_202_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_202_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14196__A1 _06057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07870__A1 _02175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_186_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13453_ _06529_ _01227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_10665_ _03991_ _04570_ _04571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_201_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_12404_ _05755_ _00952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_127_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13384_ _03663_ _06356_ _06416_ _06479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_154_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10596_ _04242_ _04507_ _04524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_103_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15123_ _00976_ net3 mod.u_cpu.rf_ram.memory\[170\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__14800__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07622__A1 _01918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12335_ _05708_ _00930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_86_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15054_ _00908_ net3 mod.u_cpu.rf_ram.memory\[192\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_141_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12266_ _05604_ _05662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_257_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14005_ _06942_ _06966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_141_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11217_ _04938_ mod.u_cpu.rf_ram.memory\[327\]\[0\] _04946_ _04947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_96_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12197_ _05588_ _05594_ _05615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_68_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09094__I _03349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07607__I _01914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14950__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_233_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11148_ _04900_ _00551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_95_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_5370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11079_ _04854_ _00528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_3_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09678__A2 _03873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09822__I _03985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14907_ _00761_ net3 mod.u_cpu.rf_ram.memory\[231\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07233__S0 _01540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_209_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11485__A2 _05130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07770__C _02077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15306__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_184_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13344__I _06121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_236_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14838_ _00692_ net3 mod.u_cpu.rf_ram.memory\[268\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_149_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_224_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3990 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_252_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_225_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_211_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14769_ _00623_ net3 mod.u_cpu.rf_ram.memory\[303\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_output6_I net6 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_205_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07310_ _01551_ _01618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_147_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10296__I0 _04313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14330__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15456__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_176_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08290_ _01882_ _02597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_189_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_220_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14187__A1 _03842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_177_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07241_ _01505_ _01544_ _01548_ _01529_ _01549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__07861__A1 _02150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12037__I1 _05468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12737__A2 _05552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07172_ mod.u_cpu.cpu.immdec.imm24_20\[3\] _01467_ _01480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09989__I0 _04091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_191_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08106__C _01830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14480__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_191_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_145_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_258_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07945__C _02252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_207_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_154_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07517__I _01743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09813_ _03768_ _03966_ _03979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_115_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_259_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_154_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09744_ _03714_ _03893_ _03926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_74_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09669__A2 _03866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09732__I _03915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09675_ _03870_ _03848_ _03871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_36_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2007 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2018 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2029 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08626_ _01486_ _02923_ _02932_ _02933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_199_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07252__I mod.u_cpu.raddr\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08557_ mod.u_cpu.rf_ram.memory\[304\]\[1\] mod.u_cpu.rf_ram.memory\[305\]\[1\] mod.u_cpu.rf_ram.memory\[306\]\[1\]
+ mod.u_cpu.rf_ram.memory\[307\]\[1\] _01994_ _02010_ _02864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_70_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_196_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07508_ _01694_ _01737_ _01738_ _01815_ _01816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_168_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_204_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08488_ _02668_ _02791_ _02794_ _02096_ _02795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_196_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10987__A1 _04238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14823__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07852__A1 _02156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07439_ _01746_ _01747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_149_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13925__A1 _06249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08083__I _01679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10450_ _04425_ _00328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_108_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11787__I0 _05311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09109_ _03385_ _03409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07604__A1 _01848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_202_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10381_ _04378_ _04379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__12534__S _05846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_191_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_12120_ _05562_ _00861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__14973__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12051_ _05498_ mod.u_cpu.rf_ram.memory\[61\]\[0\] _05516_ _05517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_123_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11002_ mod.u_cpu.rf_ram.memory\[361\]\[0\] _04658_ _04799_ _04800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_105_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15329__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10911__A1 _04172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_265_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_219_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_266_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_252_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_12953_ _06125_ _06129_ _06130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_3220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_218_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11904_ _05417_ _05401_ _05418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08258__I _02245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14353__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15479__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12884_ _06070_ mod.u_cpu.rf_ram.memory\[99\]\[1\] _06077_ _06079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_3286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07162__I _01470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07391__I0 mod.u_cpu.rf_ram.memory\[408\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_234_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_221_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14623_ _00477_ net3 mod.u_cpu.rf_ram.memory\[376\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11835_ _05366_ mod.u_cpu.rf_ram.memory\[228\]\[0\] _05368_ _05369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_2574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_199_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14554_ _00408_ net3 mod.u_cpu.rf_ram.memory\[410\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11766_ _03944_ _05322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_144_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09832__A2 _03993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1895 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14169__A1 _05780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13505_ _06561_ _01247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_159_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10717_ _04605_ _00415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_174_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_14485_ _00339_ net3 mod.u_cpu.rf_ram.memory\[445\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12508__I _05725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11697_ _05274_ _00726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_187_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_186_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13436_ _06510_ _06519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_10648_ _04559_ _00392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_173_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13392__A2 _06397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13367_ _06308_ _06463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_255_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10579_ _04506_ mod.u_cpu.rf_ram.memory\[42\]\[0\] _04512_ _04513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_142_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15106_ _00960_ net3 mod.u_cpu.rf_ram.memory\[439\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_114_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12318_ _05696_ mod.u_cpu.rf_ram.memory\[189\]\[0\] _05697_ _05698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_114_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13298_ _06289_ _06390_ _06394_ _06373_ _06395_ _06396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_108_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09348__A1 _03568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15037_ _00891_ net3 mod.u_cpu.rf_ram.memory\[1\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12249_ _05649_ _05650_ _05651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_130_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07337__I _01644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08020__A1 _02297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13783__B _06455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_228_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11950__I0 _05450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08571__A2 mod.u_cpu.rf_ram.memory\[276\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07790_ _01637_ _02098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_37_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09552__I _03773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_260_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10698__I _04578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12655__A1 _05742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_266_1313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09460_ _03388_ _03337_ _03687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_184_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08168__I _02475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_184_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_251_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08411_ _02656_ mod.u_cpu.rf_ram.memory\[446\]\[1\] _02717_ _01961_ _02718_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_240_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14846__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09391_ mod.u_arbiter.i_wb_cpu_dbus_adr\[25\] _03615_ _03628_ _03629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_184_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11523__S _05156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_205_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08342_ _02220_ _02648_ _02649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_51_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09823__A2 _03986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_220_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12418__I _05229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08273_ _02542_ _02572_ _02580_ _02491_ _02581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__07834__A1 _02110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_193_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11322__I _04995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14996__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07224_ _01531_ _01532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13758__I1 mod.u_arbiter.i_wb_cpu_rdt\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_203_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_192_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13383__A2 _03391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07155_ _01463_ _01464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_121_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_192_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14226__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08011__A1 _02316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13185__S _06126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11941__I0 _05442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_247_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14376__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08279__S _02585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07988_ mod.u_cpu.rf_ram.memory\[104\]\[0\] mod.u_cpu.rf_ram.memory\[105\]\[0\] mod.u_cpu.rf_ram.memory\[106\]\[0\]
+ mod.u_cpu.rf_ram.memory\[107\]\[0\] _02294_ _02295_ _02296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_263_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_210_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15621__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09727_ _03877_ mod.u_cpu.rf_ram.memory\[555\]\[0\] _03912_ _03913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_170_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_234_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_228_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09658_ _03857_ _03858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_43_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08078__I _01581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_216_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_188_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_70_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08609_ _02040_ _02915_ _02916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09589_ _03779_ _03786_ _03803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_230_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_208_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11620_ _05220_ _00703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_169_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_196_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11551_ _04758_ _05171_ _05175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07825__A1 _02129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_211_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15001__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_196_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10502_ _04453_ mod.u_cpu.rf_ram.memory\[442\]\[0\] _04461_ _04462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_14270_ _00124_ net3 mod.u_cpu.rf_ram.memory\[552\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_17_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11482_ _05128_ mod.u_cpu.rf_ram.memory\[286\]\[1\] _05126_ _05129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_10_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13221_ _03501_ mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat\[0\] _06327_ _06328_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_87_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10433_ _04414_ _04413_ _04415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11385__A1 _04377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13152_ mod.u_arbiter.i_wb_cpu_rdt\[27\] mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat\[11\]
+ _06263_ _06267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_109_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10364_ _04367_ _00300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_174_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__15151__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12103_ _05551_ _00855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_151_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_152_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13083_ _06205_ mod.u_cpu.rf_ram.memory\[104\]\[0\] _06224_ _06225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_10295_ _04320_ _00278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__14719__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12034_ _03728_ _04955_ _05506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_151_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08002__A1 _02293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11608__S _05211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14869__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13985_ mod.u_arbiter.i_wb_cpu_dbus_dat\[10\] _06943_ _06951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_253_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09502__A1 _03723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3050 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12936_ mod.u_cpu.cpu.genblk3.csr.timer_irq_r _06111_ _06112_ _06113_ _06063_ _06114_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XTAP_3061 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3072 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_222_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3083 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_233_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_222_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_207_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_222_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3094 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12867_ _03677_ _06066_ _06067_ _01103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_222_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11860__A2 _04378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11818_ _05357_ _00764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_14606_ _00460_ net3 mod.u_cpu.rf_ram.memory\[384\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_15586_ _01357_ net3 mod.u_arbiter.i_wb_cpu_dbus_dat\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_33_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12798_ _06022_ _01079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_14_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09805__A2 _03966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08459__I3 mod.u_cpu.rf_ram.memory\[379\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_187_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14537_ _00391_ net3 mod.u_cpu.rf_ram.memory\[41\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11749_ _03696_ _05309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_175_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14468_ _00322_ net3 mod.u_cpu.rf_ram.memory\[453\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__14249__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_179_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09569__A1 _03700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13419_ _06507_ _01215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_14399_ _00253_ net3 mod.u_cpu.rf_ram.memory\[488\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_143_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08241__A1 _02546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_192_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_154_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08960_ _03253_ _03261_ _03262_ _03264_ _03265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_88_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11128__A1 _04741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14399__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15644__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07911_ _01607_ _02215_ _02217_ _02218_ _02219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_151_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_257_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__12876__A1 _05494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08891_ _02479_ _03197_ _03198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_68_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_229_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11518__S _05153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07842_ _01741_ _02150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_96_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_245_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_216_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07773_ mod.u_cpu.rf_ram.memory\[176\]\[0\] mod.u_cpu.rf_ram.memory\[177\]\[0\] mod.u_cpu.rf_ram.memory\[178\]\[0\]
+ mod.u_cpu.rf_ram.memory\[179\]\[0\] _02048_ _02049_ _02081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_37_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09512_ _03736_ _00079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_266_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_213_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09443_ _03391_ _03674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_197_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_266_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_227_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_213_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_212_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13532__I _03292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_213_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__15024__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09374_ _03496_ mod.u_scanchain_local.module_data_in\[61\] _03613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__07530__I _01503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08325_ _01495_ _02632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_127_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08256_ _02528_ _02563_ _02564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_20_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__15174__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_193_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_192_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07207_ mod.u_cpu.raddr\[0\] _01515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08187_ _02393_ _02495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_181_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10414__I0 _04400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07138_ _01446_ _01447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_161_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13200__C _06306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08783__A2 _03089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10080_ _04162_ mod.u_cpu.rf_ram.memory\[505\]\[0\] _04165_ _04166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12867__A1 _03677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_235_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_262_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13770_ _03403_ _06771_ _03377_ _06772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_10982_ _04774_ mod.u_cpu.rf_ram.memory\[364\]\[0\] _04785_ _04786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_74_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_215_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11142__I1 mod.u_cpu.rf_ram.memory\[340\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_204_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12721_ _05588_ _05952_ _05972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_43_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_254_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_128_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_231_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15440_ _00003_ net3 mod.u_cpu.cpu.alu.add_cy_r vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_231_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12652_ _05926_ _01029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_43_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11603_ _05209_ _00697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_54_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15517__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15371_ _01146_ net3 mod.u_cpu.rf_ram.memory\[83\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_12_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12583_ _05869_ mod.u_cpu.rf_ram.memory\[157\]\[0\] _05879_ _05880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_212_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14322_ _00176_ net3 mod.u_cpu.rf_ram.memory\[526\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10653__I0 _04557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11534_ _03835_ _05164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_8_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13347__A2 _06314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14253_ _00107_ net3 mod.u_cpu.rf_ram.memory\[561\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_144_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11465_ _05116_ _00652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_184_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_256_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13204_ _06310_ _06311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_165_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14541__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10416_ _04387_ mod.u_cpu.rf_ram.memory\[456\]\[1\] _04401_ _04403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08223__A1 _02527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14184_ _01985_ _07086_ _07087_ _01400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_174_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11396_ _05070_ _00629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_124_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13135_ _06257_ _01181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_180_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_152_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10347_ _04345_ mod.u_cpu.rf_ram.memory\[467\]\[1\] _04354_ _04356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_180_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_151_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_139_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_239_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_152_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13066_ _06213_ _01156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_10278_ _04301_ _04308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11905__I0 _05413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14691__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_215_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12017_ _05494_ _05471_ _05495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09723__A1 _03711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08526__A2 _02825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_239_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08082__S0 _02171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_227_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_266_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_207_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08909__S0 _02507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15047__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12086__A2 _05388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13968_ mod.u_arbiter.i_wb_cpu_rdt\[4\] _06938_ _06928_ _03444_ _06939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_93_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_207_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09830__I _03806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_207_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12919_ _06101_ _01121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_13899_ _01453_ _06140_ _06885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13352__I _06316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_181_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15638_ _01409_ net3 mod.u_cpu.cpu.mem_bytecnt\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_222_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_221_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_222_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_210_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07350__I _01657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_210_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15197__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_194_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_194_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15569_ _01340_ net3 mod.u_arbiter.i_wb_cpu_dbus_dat\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_30_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11801__S _05344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08110_ _01592_ _02402_ _02417_ _02418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_159_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09090_ _03390_ _03391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08041_ _02058_ _02349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_163_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_266_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11349__A1 _05037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08214__A1 _02039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08181__I _01717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09962__A1 _03911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09992_ _04096_ mod.u_cpu.rf_ram.memory\[518\]\[0\] _04103_ _04104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_115_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_192_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10572__A2 _04507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_170_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08943_ mod.u_cpu.rf_ram_if.rdata0\[1\] _03248_ _01478_ _03249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_142_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12849__A1 _02523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_233_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08517__A2 _02823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08874_ mod.u_cpu.rf_ram.memory\[559\]\[1\] _03181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_215_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07525__I _01679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07825_ _02129_ mod.u_cpu.rf_ram.memory\[164\]\[0\] _02132_ _02133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_3819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_217_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07820__S0 _02125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_244_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07756_ mod.u_cpu.rf_ram.memory\[136\]\[0\] mod.u_cpu.rf_ram.memory\[137\]\[0\] mod.u_cpu.rf_ram.memory\[138\]\[0\]
+ mod.u_cpu.rf_ram.memory\[139\]\[0\] _02022_ _02063_ _02064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_53_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_198_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14414__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07687_ _01762_ _01995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_44_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_198_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09426_ _03654_ _03658_ _00072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_125_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07260__I _01497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_197_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_240_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09357_ _03598_ _03595_ _03599_ _03600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_40_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11588__A1 _04784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14564__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08308_ mod.u_cpu.rf_ram.memory\[479\]\[1\] _02615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__07256__A2 mod.u_cpu.rf_ram.memory\[478\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_205_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09288_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[10\] _03541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_100_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13329__A2 _06402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_193_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08239_ mod.u_cpu.rf_ram.memory\[525\]\[0\] _02547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_180_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_197_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11250_ _04831_ _04969_ _04970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_165_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_238_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_180_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_118_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08024__C _01916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10201_ _04245_ mod.u_cpu.rf_ram.memory\[48\]\[1\] _04252_ _04254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09953__A1 _03899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11181_ _04643_ _04922_ _04923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_122_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_121_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10132_ _04193_ mod.u_cpu.rf_ram.memory\[498\]\[0\] _04203_ _04204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_121_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13437__I _06513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_248_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14940_ _00794_ net3 mod.u_cpu.rf_ram.memory\[222\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10063_ _04140_ mod.u_cpu.rf_ram.memory\[508\]\[1\] _04152_ _04154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_209_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_212_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11512__A1 _04873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07435__I _01560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14871_ _00725_ net3 mod.u_cpu.rf_ram.memory\[251\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_75_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_169_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13822_ _06814_ _06815_ _06817_ _06820_ _06753_ _06821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_263_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12068__A2 _04845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10079__A1 _04163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12312__I0 _05692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_204_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13753_ _06726_ _06472_ _06283_ _06712_ _06757_ _06758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_1_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10796__I _03924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_189_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10965_ _04773_ _00495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_90_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12704_ _05960_ _01047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_204_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14907__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_182_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08692__A1 _02348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13684_ _06367_ _06694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_203_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10896_ _04720_ mod.u_cpu.rf_ram.memory\[378\]\[1\] _04725_ _04727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_12635_ _05914_ _01024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_15423_ _01198_ net3 mod.u_cpu.rf_ram.memory\[94\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_157_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_223_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10626__I0 _04523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15354_ _01129_ net3 mod.u_cpu.cpu.genblk3.csr.mie_mtie vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12566_ _05858_ mod.u_cpu.rf_ram.memory\[160\]\[1\] _05866_ _05868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_157_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11517_ _04732_ _05149_ _05153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_14305_ _00159_ net3 mod.u_cpu.rf_ram.memory\[535\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_102_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_129_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10237__S _04278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15285_ _00044_ net4 mod.u_scanchain_local.module_data_in\[42\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_172_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12497_ _05606_ _04309_ _05824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09097__I net5 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_176_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14236_ _00090_ net3 mod.u_cpu.rf_ram.memory\[56\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_172_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11448_ _05096_ mod.u_cpu.rf_ram.memory\[290\]\[0\] _05103_ _05104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_144_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11051__I0 _04825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08747__A2 mod.u_cpu.rf_ram.memory\[108\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13740__A2 _06425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10036__I _04133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_4_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_14167_ _07071_ _07075_ _07076_ _01393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_11379_ _04775_ _05058_ _05059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_152_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_252_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13118_ _06237_ mod.u_cpu.rf_ram.memory\[0\]\[1\] _06245_ _06247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_152_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08869__C _02518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14098_ _07028_ mod.u_cpu.rf_ram.memory\[120\]\[1\] _07030_ _07032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__13879__I0 mod.u_arbiter.i_wb_cpu_rdt\[24\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13049_ _02373_ _06201_ _06202_ _01150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_230_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_79_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_239_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14437__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_254_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_187_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07610_ _01750_ _01918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_226_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08590_ _02688_ _02895_ _02896_ _01698_ _02897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_38_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_208_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07541_ _01832_ _01849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_208_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_207_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_228_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_263_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_250_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14587__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08176__I _01745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08683__A1 _02594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07472_ mod.u_cpu.rf_ram.memory\[431\]\[0\] _01780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__07486__A2 _01793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09211_ _03478_ _00034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08109__C _02363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10490__A1 _04315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_179_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_210_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_148_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09142_ _03409_ _03436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_148_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08435__A1 _02609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12231__A2 _05637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_175_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10242__A1 _04281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09073_ _03371_ _03375_ _03376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_120_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_198_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_200_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_190_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08024_ _02329_ mod.u_cpu.rf_ram.memory\[118\]\[0\] _02331_ _01916_ _02332_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_162_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08840__S _01577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13031__I1 mod.u_cpu.rf_ram.memory\[108\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_239_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_162_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08738__A2 mod.u_cpu.rf_ram.memory\[254\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13731__A2 _06483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12362__S _05727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15212__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09735__I _03918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08779__C _02291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09975_ _03714_ _04077_ _04093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_5007 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_77_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_19 io_oeb[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_103_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_5018 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5029 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_162_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08926_ _02525_ _03229_ _03232_ _02539_ _03233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_58_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_4306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_257_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11345__I1 mod.u_cpu.rf_ram.memory\[308\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12542__I0 _05827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08857_ _02102_ _03146_ _03163_ _01739_ _03164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_57_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_218_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15362__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07808_ _01862_ _02116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_85_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2904 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08788_ mod.u_cpu.rf_ram.memory\[92\]\[1\] mod.u_cpu.rf_ram.memory\[93\]\[1\] mod.u_cpu.rf_ram.memory\[94\]\[1\]
+ mod.u_cpu.rf_ram.memory\[95\]\[1\] _01636_ _01638_ _03095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__09470__I _03695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2915 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2926 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2937 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13798__A2 _06798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07739_ _02026_ _02047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2948 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2959 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10856__I0 _04698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10750_ _04360_ _04623_ _04628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_53_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08674__A1 _02479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_240_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_201_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09409_ _03561_ _03643_ _03644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_158_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10681_ _01706_ _04581_ _04582_ _00402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_90_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12420_ _05766_ _00957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12222__A2 _05631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12351_ _05719_ _00935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_194_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12336__I _05105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13970__A2 _03614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_217_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_153_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11302_ _05006_ _00599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_154_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15070_ _00924_ net3 mod.u_cpu.rf_ram.memory\[189\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_126_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12282_ _05673_ _00912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_107_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14021_ _06942_ _06978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_11233_ mod.u_cpu.rf_ram.memory\[325\]\[1\] _04819_ _04956_ _04958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__13722__A2 _06662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09645__I _03739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_253_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08689__C _02093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11164_ _04911_ _00556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_253_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07593__C _01677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10115_ _04162_ mod.u_cpu.rf_ram.memory\[500\]\[0\] _04190_ _04191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_95_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_249_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_216_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11095_ _04457_ _04848_ _04865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_5541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__13486__B2 _03616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11336__I1 mod.u_cpu.rf_ram.memory\[30\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_209_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14923_ _00777_ net3 mod.u_cpu.rf_ram.memory\[6\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_29_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10046_ _04135_ _04142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_5574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_236_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_4851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_110_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_236_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_208_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10520__S _04473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14854_ _00708_ net3 mod.u_cpu.rf_ram.memory\[260\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_4884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4895 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13805_ _06468_ _06452_ _06779_ _06804_ _06776_ _06805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_205_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14785_ _00639_ net3 mod.u_cpu.rf_ram.memory\[295\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11997_ _05019_ _05433_ _05481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__09457__A3 _03682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_205_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_189_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13736_ _06726_ _06459_ _06741_ _06442_ _06381_ _06742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__08665__A1 _02561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07468__A2 _01775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10948_ _04762_ _00489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_260_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12461__A2 _03355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_220_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_231_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_204_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13667_ mod.u_cpu.cpu.immdec.imm19_12_20\[1\] _06678_ _06679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10879_ _04698_ mod.u_cpu.rf_ram.memory\[381\]\[1\] _04714_ _04716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_220_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_15406_ _01181_ net3 mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_176_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12618_ _05903_ _01018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13598_ mod.u_cpu.cpu.bufreg.i_sh_signed _03669_ _03693_ _06620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__10224__A1 _04230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15337_ _01112_ net3 mod.u_cpu.rf_ram.memory\[98\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12549_ _05857_ _00995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_258_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15235__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10775__A2 _04644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15268_ _00025_ net4 mod.u_arbiter.i_wb_cpu_rdt\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11024__I0 _04797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14219_ _07107_ _01416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13713__A2 _06704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15199_ _01052_ net3 mod.u_cpu.rf_ram.memory\[138\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_154_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_193_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15385__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09760_ _03747_ _03748_ _03938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_113_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_239_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09491__S _01418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08711_ mod.u_cpu.rf_ram.memory\[232\]\[1\] mod.u_cpu.rf_ram.memory\[233\]\[1\] mod.u_cpu.rf_ram.memory\[234\]\[1\]
+ mod.u_cpu.rf_ram.memory\[235\]\[1\] _01647_ _01732_ _03018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_67_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09691_ _03746_ _03710_ _03883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_94_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_255_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08642_ mod.u_cpu.rf_ram.memory\[175\]\[1\] _02949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_26_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_227_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_148_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08573_ _01949_ _02879_ _02880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_148_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_70_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_223_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07524_ _01444_ _01832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__08656__A1 _02105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08200__S0 _02507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_222_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_161_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07455_ _01762_ _01763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_161_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08408__A1 _02462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13401__A1 _06438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07386_ _01676_ _01692_ _01693_ _01694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_124_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09125_ mod.u_arbiter.i_wb_cpu_rdt\[0\] _03415_ _03422_ _03423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_194_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10066__I1 mod.u_cpu.rf_ram.memory\[507\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_198_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_198_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_148_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_191_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11963__A1 _05139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10766__A2 _04623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_198_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09056_ _03280_ _03359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_194_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_159_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09208__I0 mod.u_arbiter.i_wb_cpu_rdt\[29\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08007_ _02297_ mod.u_cpu.rf_ram.memory\[124\]\[0\] _02314_ _02315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__14602__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09465__I _03292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12763__I0 _05998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_235_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09958_ _04073_ mod.u_cpu.rf_ram.memory\[524\]\[0\] _04081_ _04082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_253_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14752__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08909_ mod.u_cpu.rf_ram.memory\[520\]\[1\] mod.u_cpu.rf_ram.memory\[521\]\[1\] mod.u_cpu.rf_ram.memory\[522\]\[1\]
+ mod.u_cpu.rf_ram.memory\[523\]\[1\] _02507_ _02543_ _03216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_213_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_218_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09889_ _03945_ _04034_ _04035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_44_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13715__I mod.u_cpu.cpu.immdec.imm19_12_20\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11920_ _05413_ mod.u_cpu.rf_ram.memory\[222\]\[0\] _05429_ _05430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_3424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07537__I3 mod.u_cpu.rf_ram.memory\[339\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12691__A2 _05319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11851_ _05364_ mod.u_cpu.rf_ram.memory\[149\]\[1\] _05378_ _05380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__15108__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_233_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11235__I _03737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10802_ _04662_ _00443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14570_ _00424_ net3 mod.u_cpu.rf_ram.memory\[402\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11782_ _05329_ mod.u_cpu.rf_ram.memory\[235\]\[1\] _05331_ _05333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_214_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08745__S _01508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_202_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_198_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13640__A1 _03297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_260_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_241_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_198_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10733_ _04608_ mod.u_cpu.rf_ram.memory\[404\]\[1\] _04614_ _04616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_13521_ _06573_ _06574_ _06575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_213_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__15258__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13452_ _03541_ _06525_ _06526_ _03547_ _06529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_185_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10664_ _04569_ _04570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07870__A2 mod.u_cpu.rf_ram.memory\[204\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12403_ _05753_ mod.u_cpu.rf_ram.memory\[176\]\[0\] _05754_ _05755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_139_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_220_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_13383_ _03665_ _03391_ _03672_ _06478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_126_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10595_ _04522_ _04523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_182_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12334_ _05696_ mod.u_cpu.rf_ram.memory\[183\]\[0\] _05707_ _05708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_15122_ _00975_ net3 mod.u_cpu.rf_ram.memory\[170\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_154_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14282__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15053_ _00907_ net3 mod.u_cpu.rf_ram.memory\[193\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_182_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12265_ _05661_ _00907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_141_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11706__A1 _04994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14004_ _06962_ _06965_ _01342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11216_ _04668_ _04945_ _04946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_12196_ _05614_ _00885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_123_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11147_ mod.u_cpu.rf_ram.memory\[33\]\[1\] _04819_ _04898_ _04900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_68_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12506__I0 _05822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11078_ _04843_ mod.u_cpu.rf_ram.memory\[350\]\[0\] _04853_ _04854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_7_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_237_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_5393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14906_ _00760_ net3 mod.u_cpu.rf_ram.memory\[231\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10029_ _03986_ _04118_ _04129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_209_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08886__A1 _02461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07233__S1 _01501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_264_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14837_ _00691_ net3 mod.u_cpu.rf_ram.memory\[26\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12809__I1 _06005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_184_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3980 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_149_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3991 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_264_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_14768_ _00622_ net3 mod.u_cpu.rf_ram.memory\[303\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__13631__A1 _06371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12434__A2 _05774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_204_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_177_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11493__I0 _05114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13719_ _06320_ _06726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_108_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_232_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13360__I _06455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14699_ _00553_ net3 mod.u_cpu.rf_ram.memory\[338\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_31_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07240_ _01545_ mod.u_cpu.rf_ram.memory\[462\]\[0\] _01547_ _01525_ _01548_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_258_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__14187__A2 _05263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07861__A2 _02153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11245__I0 _04961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_176_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14625__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_176_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07171_ mod.u_cpu.cpu.immdec.imm19_12_20\[7\] _01479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__09989__I1 mod.u_cpu.rf_ram.memory\[51\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11945__A1 _04983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_201_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_172_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13698__A1 _06421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14775__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08403__B _02709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_193_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_236_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07377__A1 _01680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09812_ _03978_ _00137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_114_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_228_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09743_ _03924_ _03925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07129__A1 _01425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12122__A1 _05563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09674_ _03778_ _03870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_223_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_215_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07533__I _01710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2008 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2019 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08625_ _02925_ _02927_ _02929_ _02931_ _02077_ _02932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_254_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08556_ _01915_ _02855_ _02862_ _01812_ _02863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15400__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_242_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_223_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07507_ _01739_ _01790_ _01814_ _01815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_168_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_211_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08487_ _01496_ mod.u_cpu.rf_ram.memory\[358\]\[1\] _02793_ _02453_ _02794_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__13270__I _06120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_211_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_196_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07438_ _01568_ _01746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_168_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_211_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07852__A2 mod.u_cpu.rf_ram.memory\[196\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_241_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13925__A2 _06901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07369_ _01550_ _01677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__15550__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_182_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09108_ _03407_ _03408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_182_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08801__A1 _02204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10380_ _03721_ _04134_ _04378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_108_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_136_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09039_ mod.u_cpu.cpu.decode.op26 _01452_ _03343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_108_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_12050_ _05515_ _03810_ _05516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_117_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07368__A1 _01658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11001_ _04527_ _04780_ _04799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__12361__A1 _05535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_81_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10911__A2 _04713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_219_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13161__I0 mod.u_arbiter.i_wb_cpu_rdt\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12952_ _06128_ _06129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08868__A1 _02455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_133_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13861__A1 _06853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07443__I _01750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11903_ _03984_ _05417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_3265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_206_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12883_ _06078_ _01108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_209_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__15080__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14622_ _00476_ net3 mod.u_cpu.rf_ram.memory\[376\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11834_ _05367_ _05335_ _05368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13613__A1 _03378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14648__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_199_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11765_ _04377_ _05320_ _05321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_53_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_14553_ _00407_ net3 mod.u_cpu.rf_ram.memory\[411\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_214_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_199_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09293__A1 _03528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15312__D _00073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1896 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10716_ _04593_ mod.u_cpu.rf_ram.memory\[407\]\[1\] _04603_ _04605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_13504_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[30\] _06557_ _06558_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[31\]
+ _06561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_11696_ _05268_ mod.u_cpu.rf_ram.memory\[254\]\[0\] _05273_ _05274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_14484_ _00338_ net3 mod.u_cpu.rf_ram.memory\[445\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_202_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13377__B1 _06458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_201_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_158_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10647_ _04557_ mod.u_cpu.rf_ram.memory\[418\]\[0\] _04558_ _04559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_13435_ _06518_ _01220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_186_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14798__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11927__A1 _05348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_220_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13366_ _06326_ _06391_ _06330_ _06462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_10578_ _04511_ _03919_ _04512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_259_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_127_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15105_ _00959_ net3 mod.u_cpu.rf_ram.memory\[174\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_155_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10245__S _04282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12317_ _05515_ _05686_ _05697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_13297_ _06301_ _06395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_127_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12727__I0 _05963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12248_ _05432_ _05650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_15036_ _00890_ net3 mod.u_cpu.rf_ram.memory\[1\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_170_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_190_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_170_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_218_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12179_ _05602_ _00880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_68_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09833__I _03994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08877__C _02083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13355__I _06450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13152__I0 mod.u_arbiter.i_wb_cpu_rdt\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_231_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08859__A1 _01471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15423__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07353__I _01660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_265_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10666__A1 _04542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_236_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08410_ _01709_ _02716_ _02717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_252_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09390_ _03564_ _03625_ _03627_ _03628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_197_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_224_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_205_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08341_ mod.u_cpu.rf_ram.memory\[511\]\[1\] _02648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__10418__A1 _03942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11466__I0 _05108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_178_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15573__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09284__A1 mod.u_cpu.cpu.ctrl.o_ibus_adr\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08272_ _02545_ _02575_ _02579_ _02555_ _02580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_193_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07223_ mod.u_cpu.raddr\[3\] _01531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_165_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13907__A2 _06661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10219__I _04176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_177_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11769__I1 _05230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07154_ _01462_ _01463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__13383__A3 _03672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07956__C _01766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_195_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08634__I1 mod.u_cpu.rf_ram.memory\[189\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07988__I3 mod.u_cpu.rf_ram.memory\[107\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_145_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12718__I0 _05966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07528__I _01677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_236_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12370__S _05733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09743__I _03924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_259_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07987_ _01854_ _02295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_75_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13143__I0 mod.u_arbiter.i_wb_cpu_rdt\[23\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_170_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_256_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09726_ _03902_ _03911_ _03912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08359__I _01762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09898__I0 _04036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13843__A1 _06677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10657__A1 _04290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_255_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09657_ _03856_ _03848_ _03857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08608_ mod.u_cpu.rf_ram.memory\[128\]\[1\] mod.u_cpu.rf_ram.memory\[129\]\[1\] mod.u_cpu.rf_ram.memory\[130\]\[1\]
+ mod.u_cpu.rf_ram.memory\[131\]\[1\] _02638_ _02067_ _02915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_09588_ _03739_ _03802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_43_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_247_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_187_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08539_ _01843_ _02845_ _02846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_196_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11550_ _05174_ _00679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_168_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11082__A1 _04808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_184_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_196_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14940__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10501_ _04322_ _04443_ _04461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11481_ _05107_ _05128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_156_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10129__I _03858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_183_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13220_ _06122_ _06123_ _06327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_137_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10432_ _03898_ _04414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_183_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11385__A2 _05062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__12582__A1 _05515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_178_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13151_ _06266_ _01188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_10363_ _04365_ mod.u_cpu.rf_ram.memory\[464\]\[0\] _04366_ _04367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_124_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12102_ _05550_ mod.u_cpu.rf_ram.memory\[67\]\[1\] _05547_ _05551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07438__I _01568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13082_ _03932_ _06223_ _06224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10294_ _04298_ mod.u_cpu.rf_ram.memory\[475\]\[0\] _04319_ _04320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_215_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08978__B mod.u_cpu.cpu.state.init_done vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12033_ _05505_ _00831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_78_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_266_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08002__A2 _02296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14320__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15446__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_265_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13134__I0 mod.u_arbiter.i_wb_cpu_rdt\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13175__I _06281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07761__A1 _02046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13834__A1 _06651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13984_ _06949_ _06950_ _01337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_46_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_247_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_218_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09502__A2 _03727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3040 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11696__I0 _05268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3051 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14470__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12935_ _01434_ _06113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__15596__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3062 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3073 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3084 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_234_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3095 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_234_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12866_ mod.u_cpu.cpu.state.ibus_cyc _06066_ _06046_ _06067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_206_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07901__I _02091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_248_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11448__I0 _05096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14605_ _00459_ net3 mod.u_cpu.rf_ram.memory\[385\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11817_ _05342_ mod.u_cpu.rf_ram.memory\[230\]\[0\] _05356_ _05357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_159_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15585_ _01356_ net3 mod.u_arbiter.i_wb_cpu_dbus_dat\[27\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09266__A1 _03506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12797_ _06010_ mod.u_cpu.rf_ram.memory\[12\]\[0\] _06021_ _06022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_1671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14536_ _00390_ net3 mod.u_cpu.rf_ram.memory\[41\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_261_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11748_ _05308_ _00743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_144_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10039__I _04136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09018__A1 _03259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14467_ _00321_ net3 mod.u_cpu.rf_ram.memory\[454\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11679_ _05261_ _00721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_174_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_13418_ _06351_ mod.u_cpu.rf_ram.memory\[339\]\[0\] _06506_ _06507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_14398_ _00252_ net3 mod.u_cpu.rf_ram.memory\[488\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_155_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13349_ _06422_ _06445_ _06446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_66_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13794__B _06486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15019_ _00873_ net3 mod.u_cpu.rf_ram.memory\[206\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_07910_ _01746_ _02218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_08890_ mod.u_cpu.rf_ram.memory\[565\]\[1\] _03197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_97_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12876__A2 _05263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_190_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07841_ _01488_ _02149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_111_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14813__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_238_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07772_ _01661_ _02080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08179__I _02010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09511_ mod.u_cpu.rf_ram.memory\[9\]\[1\] _03735_ _03729_ _03736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_65_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_266_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_237_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_225_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09442_ _03663_ _03666_ _03669_ _03672_ _03673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_37_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_240_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_253_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__14963__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09373_ _03489_ _03611_ _03612_ _00065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_40_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08324_ _02347_ _02631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_178_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10111__I0 _04178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_221_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_193_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_177_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15319__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09009__A1 _01430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08255_ mod.u_cpu.rf_ram.memory\[533\]\[0\] _02563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_220_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_197_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12365__S _05727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08480__A2 _02779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07206_ _01508_ mod.u_cpu.rf_ram.memory\[452\]\[0\] _01513_ _01514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_181_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08186_ _01705_ _02494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_165_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10414__I1 mod.u_cpu.rf_ram.memory\[456\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07137_ _01445_ _01446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_146_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14343__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__15469__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10178__I0 _04215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09473__I _03698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_247_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14069__A1 mod.u_arbiter.i_wb_cpu_rdt\[31\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14493__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_181_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11508__I _05107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13116__I0 _06230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_263_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08310__C _01751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10412__I _04347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_261_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_229_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11678__I0 _05250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09709_ _03898_ _03899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_216_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10981_ _04784_ _04759_ _04785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_90_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09496__A1 _03718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_216_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_245_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12720_ _03698_ _05971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_216_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_204_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10350__I0 _04348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_230_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_188_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12651_ _05918_ mod.u_cpu.rf_ram.memory\[146\]\[0\] _05925_ _05926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_247_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_180_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11243__I _03967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_208_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11602_ _05208_ mod.u_cpu.rf_ram.memory\[266\]\[1\] _05206_ _05209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_145_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10102__I0 _04162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12582_ _05515_ _05374_ _05879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_15370_ _01145_ net3 mod.u_cpu.rf_ram.memory\[108\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_141_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09263__A4 _03498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14321_ _00175_ net3 mod.u_cpu.rf_ram.memory\[527\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11533_ _05163_ _00673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_168_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09648__I _03849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11464_ _05114_ mod.u_cpu.rf_ram.memory\[288\]\[0\] _05115_ _05116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_14252_ _00106_ net3 mod.u_cpu.rf_ram.memory\[561\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_99_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_13203_ _06118_ _06309_ _06310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_10415_ _04402_ _00316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11602__I0 _05208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14183_ _07026_ _07086_ _07087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_11395_ _05069_ mod.u_cpu.rf_ram.memory\[300\]\[1\] _05067_ _05070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_139_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13134_ mod.u_arbiter.i_wb_cpu_rdt\[19\] mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat\[3\]
+ _06253_ _06257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_48_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10346_ _04355_ _00294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_3_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14836__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07982__A1 _02283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_174_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13065_ _06205_ mod.u_cpu.rf_ram.memory\[106\]\[0\] _06212_ _06213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_65_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10277_ _03769_ _04307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_12016_ _03827_ _05494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_79_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_266_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09723__A2 _03788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08082__S1 _02267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_239_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_266_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_253_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__14986__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__08909__S1 _02543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13967_ _06937_ _06938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_222_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12918_ mod.u_cpu.rf_ram.memory\[389\]\[1\] _06005_ _06099_ _06101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_94_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_235_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_13898_ _01435_ _06881_ _06847_ _01317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_73_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_222_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15637_ _01408_ net3 mod.u_cpu.cpu.state.o_cnt\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12849_ _02523_ _03742_ _06054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_34_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_210_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_203_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15568_ _01339_ net3 mod.u_arbiter.i_wb_cpu_dbus_dat\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_175_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10992__I _03917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14519_ _00373_ net3 mod.u_cpu.rf_ram.memory\[428\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_202_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_147_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15499_ _01270_ net3 mod.u_arbiter.i_wb_cpu_dbus_adr\[19\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__14366__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08040_ _02347_ _02348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_266_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_200_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13301__C _06398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15611__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09411__A1 mod.u_arbiter.i_wb_cpu_dbus_adr\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08845__S0 _02349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_192_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09991_ _03951_ _04087_ _04103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_116_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07973__A1 _02079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_192_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08942_ _03247_ mod.u_cpu.rf_ram.regzero _03248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__12712__I _05937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_229_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08873_ _02478_ mod.u_cpu.rf_ram.memory\[556\]\[1\] _03179_ _03180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_96_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_218_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07725__A1 _01992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_245_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07824_ _02130_ _02131_ _02132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_3809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07820__S1 _02127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07755_ _01960_ _02063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09478__A1 _01660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_231_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07686_ _01993_ _01994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_241_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_213_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_212_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07541__I _01832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07584__S0 _01843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15141__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09425_ mod.u_arbiter.i_wb_cpu_dbus_adr\[30\] _03561_ _03656_ _03657_ _03409_ _03658_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_198_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_198_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14709__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13699__B _06707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09356_ _03598_ _03586_ _03594_ _03599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_200_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11588__A2 _05191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08307_ _02566_ mod.u_cpu.rf_ram.memory\[476\]\[1\] _02613_ _02614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_21_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09287_ _03528_ _03539_ _03540_ _00049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_139_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10608__S _04529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_176_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08238_ _02477_ _02546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_138_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15291__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_176_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14859__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12537__A1 _05642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_193_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08169_ _02047_ _02477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_119_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_88_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08836__S0 _02421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_180_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10200_ _04253_ _00250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_107_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11180_ _04379_ _04779_ _04922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_122_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10131_ _04201_ _04202_ _04203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_216_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10062_ _04153_ _00212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11899__I0 _05413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_197_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07716__A1 _01729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14870_ _00724_ net3 mod.u_cpu.rf_ram.memory\[251\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_76_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_248_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_235_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_217_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14239__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13821_ _06818_ _06819_ _06332_ _06820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_63_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11276__A1 _03755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_204_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13752_ _06666_ _06671_ _06756_ _06757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_141_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_217_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10964_ _04772_ mod.u_cpu.rf_ram.memory\[367\]\[1\] _04770_ _04773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_216_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07451__I _01758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_182_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_44_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_231_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_188_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12703_ mod.u_cpu.rf_ram.memory\[13\]\[0\] _05622_ _05959_ _05960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_44_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_204_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13683_ _06482_ _06475_ _06693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08692__A2 _02998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10895_ _04726_ _00472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__14389__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_188_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11028__A1 _04817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15422_ _01197_ net3 mod.u_cpu.cpu.bufreg.i_sh_signed vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_54_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12634_ _05907_ mod.u_cpu.rf_ram.memory\[14\]\[1\] _05912_ _05914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_54_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15634__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12776__A1 _03960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10626__I1 mod.u_cpu.rf_ram.memory\[422\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15353_ _01128_ net3 mod.u_cpu.cpu.genblk3.csr.mstatus_mie vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_180_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12565_ _05867_ _01001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_184_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14304_ _00158_ net3 mod.u_cpu.rf_ram.memory\[535\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_106_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11516_ _05152_ _00667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_141_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15284_ _00043_ net4 mod.u_scanchain_local.module_data_in\[41\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_106_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12496_ _05823_ _00976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_171_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12528__A1 _01574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13829__S _06335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13576__I0 mod.u_arbiter.i_wb_cpu_dbus_adr\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14235_ _00089_ net3 mod.u_cpu.rf_ram.memory\[570\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10317__I _04308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11447_ _04831_ _05089_ _05103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_171_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11378_ _04995_ _05058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_14166_ _06046_ _07076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13740__A3 _06458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07955__A1 _02249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_217_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__13628__I _06640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13117_ _06246_ _01174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_10329_ _04326_ mod.u_cpu.rf_ram.memory\[46\]\[0\] _04342_ _04343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_124_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_258_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15014__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14097_ _07031_ _01369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_112_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07626__I _01710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13879__I1 mod.u_arbiter.i_wb_cpu_rdt\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13048_ _06032_ _06201_ _06202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_39_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_152_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_266_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_227_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09841__I _03915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15164__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_208_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_14999_ _00853_ net3 mod.u_cpu.rf_ram.memory\[66\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__13363__I _06458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07540_ _01457_ _01848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08457__I _01660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_223_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08132__A1 _01819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07361__I _01491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_223_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07471_ _01778_ _01779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_35_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14205__A1 _07076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08683__A2 _02986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_210_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09210_ mod.u_arbiter.i_wb_cpu_rdt\[30\] mod.u_arbiter.i_wb_cpu_dbus_dat\[27\] _03474_
+ _03478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_50_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_72_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_37_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09141_ _03409_ _03435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_148_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12707__I _05694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09632__A1 _03834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08192__I _02216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10242__A2 _04263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09072_ _03374_ _03375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_198_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08125__C _02415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08023_ _01863_ _02330_ _02331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_135_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_239_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07946__A1 _02174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09974_ _04092_ _00185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_170_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5008 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07536__I _01503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5019 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08925_ _02533_ mod.u_cpu.rf_ram.memory\[542\]\[1\] _03231_ _02537_ _03232_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_170_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_4307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11058__I _03984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15507__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08856_ _03151_ _03153_ _03162_ _01891_ _03163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_58_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_217_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08371__A1 _02665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08795__C _02660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07807_ _01635_ _02115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_3639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2905 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08787_ _01662_ _03093_ _03094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2916 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2927 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_260_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07738_ _01890_ _02046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_2938 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14531__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2949 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08123__A1 _02411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_213_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08674__A2 mod.u_cpu.rf_ram.memory\[212\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07669_ _01484_ _01977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_81_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_214_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_197_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09408_ _03642_ _03638_ _03643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_186_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10680_ _04542_ _04581_ _04582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_213_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_198_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_201_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14681__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_199_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09339_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[17\] mod.u_cpu.cpu.ctrl.o_ibus_adr\[16\] mod.u_cpu.cpu.ctrl.o_ibus_adr\[15\]
+ mod.u_cpu.cpu.ctrl.o_ibus_adr\[14\] _03585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XANTENNA__10608__I1 _04532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_205_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08316__B _02622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_205_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_138_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12350_ _05711_ mod.u_cpu.rf_ram.memory\[181\]\[1\] _05717_ _05719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_193_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11301_ _04999_ mod.u_cpu.rf_ram.memory\[315\]\[1\] _05004_ _05006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__13707__B1 _06493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13558__I0 mod.u_arbiter.i_wb_cpu_dbus_adr\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12281_ _05662_ mod.u_cpu.rf_ram.memory\[190\]\[0\] _05672_ _05673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_112_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15037__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11232_ _04957_ _00578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13183__A1 _03500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14020_ _06975_ _06977_ _01346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_175_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12352__I _05629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11163_ _04901_ mod.u_cpu.rf_ram.memory\[336\]\[0\] _04910_ _04911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_136_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10792__I0 _04637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10114_ _04189_ _04164_ _04190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11094_ _04802_ _04864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__15187__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_88_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14922_ _00776_ net3 mod.u_cpu.rf_ram.memory\[6\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10045_ _04141_ _00207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_88_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_264_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10801__S _04659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_212_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_152_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14853_ _00707_ net3 mod.u_cpu.rf_ram.memory\[261\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_4874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_263_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15315__D mod.u_cpu.rf_ram_if.wdata1_r\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4896 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13804_ _06803_ _06714_ _06804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_217_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_205_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14784_ _00638_ net3 mod.u_cpu.rf_ram.memory\[295\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11996_ _05480_ _00819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_189_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09162__I0 _03449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12997__A1 _06166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13735_ _06739_ _03424_ _06740_ _06741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_45_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12997__B2 _05780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_204_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10947_ _04756_ mod.u_cpu.rf_ram.memory\[370\]\[1\] _04760_ _04762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_205_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__12461__A3 _05798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_205_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_204_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_204_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13666_ _06415_ _06678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_143_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10878_ _01859_ _04714_ _04715_ _00466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__12749__A1 _05843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_176_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_223_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15405_ _01180_ net3 mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_12617_ _05891_ mod.u_cpu.rf_ram.memory\[152\]\[1\] _05901_ _05903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XPHY_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__09614__A1 _03767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_13597_ _03659_ _03694_ _06619_ _01281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_185_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10224__A2 _04269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15336_ _01111_ net3 mod.u_cpu.rf_ram.memory\[89\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12548_ _05855_ mod.u_cpu.rf_ram.memory\[163\]\[0\] _05856_ _05857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_185_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10047__I _04142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15267_ _00024_ net4 mod.u_arbiter.i_wb_cpu_rdt\[22\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_172_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12479_ _05694_ _05812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__14210__I1 _06221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14218_ _03699_ mod.u_cpu.rf_ram.memory\[249\]\[0\] _07106_ _07107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__11024__I1 mod.u_cpu.rf_ram.memory\[358\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15198_ _01051_ net3 mod.u_cpu.rf_ram.memory\[138\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07928__A1 _02175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14404__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14149_ _03822_ _05254_ _07064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_67_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_259_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_230_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08710_ _01991_ _03017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_6_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11488__A1 _05133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09690_ _03882_ _00111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__14554__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_254_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08641_ _02111_ mod.u_cpu.rf_ram.memory\[172\]\[1\] _02947_ _02948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_265_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08187__I _02393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10510__I _04429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_242_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08572_ mod.u_cpu.rf_ram.memory\[279\]\[1\] _02879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_187_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08105__A1 _02411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_82_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_228_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07523_ mod.u_cpu.rf_ram.memory\[344\]\[0\] mod.u_cpu.rf_ram.memory\[345\]\[0\] mod.u_cpu.rf_ram.memory\[346\]\[0\]
+ mod.u_cpu.rf_ram.memory\[347\]\[0\] _01826_ _01830_ _01831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__08200__S1 _02473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_211_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07454_ _01700_ _01762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_62_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_211_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_210_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_179_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_210_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07385_ _01445_ _01693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_176_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08408__A2 mod.u_cpu.rf_ram.memory\[444\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13401__A2 _06493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_210_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09124_ _03392_ _03420_ _03421_ _03422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_202_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09081__A2 _03378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_191_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11963__A2 _03996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09055_ _03354_ _03357_ _03358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_191_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_191_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_163_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08006_ _02298_ _02313_ _02314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_144_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07919__A1 _02070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_103_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_249_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09957_ _03905_ _04062_ _04081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_104_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_213_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08908_ _02449_ _03207_ _03214_ _02469_ _03215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_103_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09888_ _03823_ _04033_ _04034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07147__A2 _01451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08344__A1 _02597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08839_ _03142_ _03143_ _03144_ _03145_ _02391_ _01552_ _03146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_3425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_245_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08097__I _02154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11850_ _05379_ _00774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_261_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_199_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12979__A1 _01453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10801_ mod.u_cpu.rf_ram.memory\[393\]\[1\] _04661_ _04659_ _04662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_2757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_198_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__10829__I1 mod.u_cpu.rf_ram.memory\[388\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11781_ _05332_ _00752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09844__A1 _03752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12548__S _05856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_202_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13640__A2 _03681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_198_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_198_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13520_ mod.u_arbiter.i_wb_cpu_dbus_adr\[2\] _03669_ _06574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10732_ _04615_ _00420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_242_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_198_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_158_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13451_ _06528_ _01226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_10663_ _04568_ _04569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_220_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_185_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_167_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12402_ _05300_ _05726_ _05754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11403__A1 _04792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13382_ _06457_ _06460_ _06477_ _01208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_142_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10594_ _04247_ _04522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_182_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__14427__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15121_ _00974_ net3 mod.u_cpu.rf_ram.memory\[171\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_154_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12333_ _03879_ _05703_ _05707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_108_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15052_ _00906_ net3 mod.u_cpu.rf_ram.memory\[193\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_108_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12264_ _05660_ mod.u_cpu.rf_ram.memory\[193\]\[1\] _05658_ _05661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_99_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_181_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13178__I _06284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11706__A2 _05279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14003_ mod.u_arbiter.i_wb_cpu_rdt\[13\] _06964_ _06958_ mod.u_arbiter.i_wb_cpu_dbus_dat\[13\]
+ _06965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_123_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_218_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11215_ _04905_ _04945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_253_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12195_ _05609_ mod.u_cpu.rf_ram.memory\[202\]\[1\] _05612_ _05614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__14577__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08583__A1 _01722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07386__A2 _01692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11146_ _04899_ _00550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_68_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_150_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_89_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11077_ _04852_ _04848_ _04853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_153_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_7_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_209_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10517__I0 _04467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_209_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08335__A1 _02597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07904__I _01701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_236_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_14905_ _00759_ net3 mod.u_cpu.rf_ram.memory\[232\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_49_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10028_ _04128_ _00203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_5394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_49_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10142__A1 _04209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11190__I0 _04916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08886__A2 mod.u_cpu.rf_ram.memory\[574\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14836_ _00690_ net3 mod.u_cpu.rf_ram.memory\[26\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_4693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3970 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3981 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_229_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3992 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_251_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_14767_ _00621_ net3 mod.u_cpu.rf_ram.memory\[304\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_189_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11979_ _05469_ _00813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09835__A1 _03991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11642__A1 _05110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13718_ _06723_ _06123_ _06724_ _06725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__15202__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11493__I1 mod.u_cpu.rf_ram.memory\[284\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_177_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_220_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14698_ _00552_ net3 mod.u_cpu.rf_ram.memory\[338\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_177_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_220_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_220_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13649_ _06404_ _06661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_176_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07170_ _01449_ _01478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_192_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_118_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_258_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11945__A2 _03837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15352__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15319_ _01098_ net3 mod.u_cpu.raddr\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07795__B _02102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_184_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08403__C _02606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10756__I0 _04622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08574__A1 _01697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07377__A2 _01684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09811_ _03964_ mod.u_cpu.rf_ram.memory\[546\]\[1\] _03976_ _03978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_140_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12720__I _03698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09742_ _03923_ _03924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10508__I0 _04453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_228_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07814__I _01719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12122__A2 _03843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_255_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09673_ _03869_ _00107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_67_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_227_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13870__A2 _06862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2009 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08624_ _02074_ _02930_ _01602_ _02931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_94_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_243_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08555_ _01981_ _02858_ _02861_ _01929_ _02862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_78_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13551__I _06583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_211_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07506_ _01791_ _01800_ _01813_ _01814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_08486_ _02672_ _02792_ _02793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_243_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_223_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_196_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_167_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_243_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_196_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07437_ _01744_ _01745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_51_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_210_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_206_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_202_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_202_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07368_ _01658_ _01668_ _01675_ _01676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_136_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09107_ _03405_ _03406_ _03407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_136_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07299_ _01539_ _01607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__08801__A2 mod.u_cpu.rf_ram.memory\[68\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09476__I _03701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_184_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_163_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08380__I _02591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09038_ mod.u_cpu.cpu.decode.op22 _03342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_124_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08565__A1 _01956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_250_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11000_ _04798_ _00505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12361__A2 _05726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_266_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_219_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_218_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__13310__A1 _06403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13161__I1 mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12951_ _06126_ _03424_ _06127_ _06128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_3211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11172__I0 _04916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11902_ _05416_ _00789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_206_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__15225__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_248_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12882_ _06073_ mod.u_cpu.rf_ram.memory\[99\]\[0\] _06077_ _06078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_3266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14621_ _00475_ net3 mod.u_cpu.rf_ram.memory\[377\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11833_ _03959_ _05367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_2554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_233_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11182__S _04923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_260_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_198_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14552_ _00406_ net3 mod.u_cpu.rf_ram.memory\[411\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11764_ _04227_ _05319_ _05320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_1864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_202_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_202_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13503_ _06560_ _01246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_159_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15375__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1897 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10715_ _01730_ _04603_ _04604_ _00414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_187_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14483_ _00337_ net3 mod.u_cpu.rf_ram.memory\[446\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11695_ _04852_ _05255_ _05273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_186_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13377__A1 _06471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13377__B2 _06395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13434_ _03507_ _06511_ _06514_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[4\] _06518_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_139_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10646_ _04281_ _04534_ _04558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_167_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11927__A2 _05434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_259_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13365_ _03664_ _03663_ _06356_ _06461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_10_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10577_ _04250_ _04511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_155_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_15104_ _00958_ net3 mod.u_cpu.rf_ram.memory\[174\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_182_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08290__I _01882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12316_ _05695_ _05696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_115_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13296_ _06313_ _06393_ _06389_ _06394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_6_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15035_ _00889_ net3 mod.u_cpu.rf_ram.memory\[200\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_114_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12247_ _03967_ _05649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_123_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10738__I0 _04608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_190_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_122_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12178_ _05575_ mod.u_cpu.rf_ram.memory\[204\]\[0\] _05601_ _05602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_151_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13636__I _06412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11129_ _04883_ mod.u_cpu.rf_ram.memory\[342\]\[0\] _04888_ _04889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_116_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_237_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_209_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11163__I0 _04901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11156__I _04905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13572__S _06604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_264_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__11863__A1 _05355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08666__S _02294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10666__A2 _04571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_266_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_4490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14101__I0 _07021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14819_ _00673_ net3 mod.u_cpu.rf_ram.memory\[278\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07382__I2 mod.u_cpu.rf_ram.memory\[398\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11092__S _04860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10418__A2 _04335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08340_ _02559_ mod.u_cpu.rf_ram.memory\[508\]\[1\] _02646_ _02647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__12663__I0 _05923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08271_ _02550_ mod.u_cpu.rf_ram.memory\[542\]\[0\] _02577_ _02578_ _02579_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_33_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_225_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_192_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07222_ _01505_ _01514_ _01526_ _01529_ _01530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__14742__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09036__A2 _03259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_203_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07153_ _01461_ _01462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_157_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_199_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_146_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08795__A1 _02465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_195_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14892__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08133__C _01828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12718__I1 mod.u_cpu.rf_ram.memory\[138\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10235__I _03968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_195_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_160_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_154_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_141_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10171__S _04229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15248__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07986_ _01864_ _02294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_68_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09725_ _03910_ _03911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_228_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_210_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09656_ _03744_ _03856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10657__A2 _04437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_167_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14272__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08607_ _01481_ _02758_ _02913_ _01469_ _02914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_43_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12098__S _05547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_215_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__15398__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09587_ _03801_ _00089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_231_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_203_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_242_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_179_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08538_ mod.u_cpu.rf_ram.memory\[293\]\[1\] _02845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_151_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_196_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11082__A2 _03975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08469_ _01852_ _02768_ _02775_ _01887_ _02776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_10_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_259_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_211_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_196_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10500_ _04460_ _00343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_11480_ _05127_ _00656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_149_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11909__A2 _05371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10431_ _04412_ _04380_ _04413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_137_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_192_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07719__I _02026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13150_ mod.u_arbiter.i_wb_cpu_rdt\[26\] mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat\[10\]
+ _06263_ _06266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_152_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12582__A2 _05374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10362_ _04209_ _04353_ _04366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_109_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_191_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12101_ _05549_ _05550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_191_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13081_ _05630_ _06223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_10293_ _03791_ _04303_ _04319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_5_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_254_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09586__I0 _03800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12032_ _05501_ mod.u_cpu.rf_ram.memory\[19\]\[1\] _05503_ _05505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_151_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13456__I _06510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_266_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12360__I _05725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07454__I _01700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_266_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_219_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13134__I1 mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07761__A2 _02068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13983_ mod.u_arbiter.i_wb_cpu_rdt\[8\] _06938_ _06947_ mod.u_arbiter.i_wb_cpu_dbus_dat\[8\]
+ _06950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_93_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14615__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_265_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13834__A2 _06829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11905__S _05418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_207_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3030 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12934_ mod.u_cpu.cpu.genblk3.csr.mie_mtie mod.u_cpu.cpu.genblk3.csr.mstatus_mie
+ mod.timer_irq _06112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__11696__I1 mod.u_cpu.rf_ram.memory\[254\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3041 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12893__I0 _06073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3052 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_262_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3063 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3074 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3085 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12865_ _06063_ _06065_ _06066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_3096 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14604_ _00458_ net3 mod.u_cpu.rf_ram.memory\[385\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__13598__A1 mod.u_cpu.cpu.bufreg.i_sh_signed vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11816_ _05355_ _05335_ _05356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__08285__I _02591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_261_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14765__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15584_ _01355_ net3 mod.u_arbiter.i_wb_cpu_dbus_dat\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12645__I0 _05918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_199_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12796_ _05870_ _03905_ _06021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_199_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_226_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_199_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14535_ _00389_ net3 mod.u_cpu.rf_ram.memory\[420\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11747_ _05304_ mod.u_cpu.rf_ram.memory\[23\]\[1\] _05306_ _05308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_1694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_175_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_230_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_202_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14466_ _00320_ net3 mod.u_cpu.rf_ram.memory\[454\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_31_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11678_ _05250_ mod.u_cpu.rf_ram.memory\[256\]\[1\] _05259_ _05261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_175_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13417_ _05732_ _04847_ _06506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10256__S _04291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10629_ _04547_ _00385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13070__I0 _06205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14397_ _00251_ net3 mod.u_cpu.rf_ram.memory\[48\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_183_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08777__A1 _02329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13770__A1 _03403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13348_ _06433_ _06440_ _06444_ _06401_ _06445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_143_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10584__A1 _04233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13279_ _06116_ _06377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_170_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08529__A1 _02148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15018_ _00872_ net3 mod.u_cpu.rf_ram.memory\[206\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09577__I0 _03764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08888__C _02505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_69_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_155_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07840_ _01482_ _02148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_69_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07364__I _01671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14295__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_231_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07771_ _02039_ _02062_ _02078_ _02079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__11136__I0 _04880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15540__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09510_ _03734_ _03735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_265_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12884__I0 _06070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08701__A1 _02063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09441_ _03670_ _03403_ _03671_ _03252_ _03672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_52_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_252_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_266_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_225_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_224_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09372_ _03563_ mod.u_scanchain_local.module_data_in\[60\] _03517_ mod.u_arbiter.i_wb_cpu_dbus_adr\[23\]
+ _03612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_36_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_240_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08323_ _02039_ _02608_ _02629_ _02630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_149_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_166_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08254_ mod.u_cpu.rf_ram.memory\[528\]\[0\] mod.u_cpu.rf_ram.memory\[529\]\[0\] mod.u_cpu.rf_ram.memory\[530\]\[0\]
+ mod.u_cpu.rf_ram.memory\[531\]\[0\] _02560_ _02561_ _02562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_123_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07967__C _02252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_177_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_193_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07205_ _01511_ _01512_ _01513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08185_ _02470_ _02492_ _01447_ _02493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_146_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_229_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_174_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08768__A1 _02316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_174_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13761__A1 _03686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07136_ _01444_ _01445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_106_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_165_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15070__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14638__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13276__I _06300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_248_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14069__A2 _06940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07274__I _01581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07969_ _01742_ _02268_ _02276_ _02207_ _02277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_247_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_228_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09708_ _03697_ _03898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_216_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11827__A1 _05348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14101__S _07033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_210_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14788__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10980_ _03903_ _04784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09496__A2 _03721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_244_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_249_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_216_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09639_ _03842_ _03843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_167_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_231_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_216_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_243_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12650_ _05293_ _05920_ _05925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12627__I0 _05904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11601_ _05177_ _05208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_19_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12581_ _05878_ _01006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_169_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10102__I1 mod.u_cpu.rf_ram.memory\[502\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_230_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11460__S _05111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14320_ _00174_ net3 mod.u_cpu.rf_ram.memory\[527\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11532_ _05162_ mod.u_cpu.rf_ram.memory\[278\]\[1\] _05160_ _05163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_168_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_183_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_168_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14251_ _00105_ net3 mod.u_cpu.rf_ram.memory\[562\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12004__A1 _03834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11463_ _04838_ _04996_ _05115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_109_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_221_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13202_ _06308_ _06309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_139_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08759__A1 _02352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08303__S0 _02593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07449__I _01515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15413__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10414_ _04400_ mod.u_cpu.rf_ram.memory\[456\]\[0\] _04401_ _04402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_109_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14182_ _03822_ _05124_ _07086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_165_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11394_ _05031_ _05069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_178_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10566__A1 _04439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_174_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_256_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_124_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13133_ _06256_ _01180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_139_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10345_ _04348_ mod.u_cpu.rf_ram.memory\[467\]\[0\] _04354_ _04355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_99_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13064_ _03918_ _06092_ _06212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10276_ _04306_ _00273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10318__A1 _04172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11366__I0 _05050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13186__I _06292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_151_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15563__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12015_ _05493_ _00825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_79_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_266_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07184__I _01491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08931__A1 _02546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11118__I0 _04880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_219_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_207_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_247_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13966_ _05801_ _06937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_98_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_207_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_111_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_207_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12917_ _06100_ _01120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12491__A1 _05334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_234_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13897_ _03342_ _06881_ _06856_ _01316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_206_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12848_ _06052_ _06053_ _01098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_61_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15636_ _01407_ net3 mod.u_cpu.cpu.state.o_cnt_r\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_22_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15567_ _01338_ net3 mod.u_arbiter.i_wb_cpu_dbus_dat\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_226_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12779_ _05998_ mod.u_cpu.rf_ram.memory\[132\]\[1\] _06007_ _06009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_261_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_203_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13991__A1 _03449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14518_ _00372_ net3 mod.u_cpu.rf_ram.memory\[428\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_175_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15498_ _01269_ net3 mod.u_arbiter.i_wb_cpu_dbus_adr\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_159_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14449_ _00303_ net3 mod.u_cpu.rf_ram.memory\[463\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_174_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15093__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13594__I1 mod.u_arbiter.i_wb_cpu_dbus_adr\[30\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09411__A2 _03561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08845__S1 _02393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_1245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09990_ _04102_ _00191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_116_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08941_ mod.u_cpu.rf_ram.rdata\[0\] _03247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_131_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_237_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11357__I0 _05032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08411__C _01961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08872_ _02479_ _03178_ _03179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07308__B _01613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14930__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07725__A2 _02021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08922__A1 _02527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07823_ mod.u_cpu.rf_ram.memory\[165\]\[0\] _02131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_96_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_229_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_38_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07754_ _02045_ _02052_ _02056_ _02061_ _01818_ _02062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_226_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07822__I _01744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07489__A1 _01779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07685_ _01645_ _01993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_64_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_253_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07584__S1 _01838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09424_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[30\] _03648_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[28\]
+ _03637_ _03657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_225_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_213_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_213_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_205_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_241_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12234__A1 _03727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09355_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[20\] _03598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_100_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_212_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14310__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08306_ _02593_ _02612_ _02613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_127_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15436__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09286_ _03535_ mod.u_scanchain_local.module_data_in\[46\] _03536_ mod.u_arbiter.i_wb_cpu_dbus_adr\[9\]
+ _03540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_165_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_197_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09650__A2 _03851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08237_ _02325_ _02545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_14_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_197_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12537__A2 _05849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_197_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13585__I1 mod.u_arbiter.i_wb_cpu_dbus_adr\[26\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08168_ _02475_ _02476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_147_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11596__I0 _05194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_180_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14460__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10399__I1 _04383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08836__S1 _02393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15586__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07413__A1 _01696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07119_ mod.u_cpu.cpu.decode.co_mem_word _01428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08099_ mod.u_cpu.rf_ram.memory\[21\]\[0\] _02407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_49_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_192_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_171_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10130_ _04142_ _04202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_238_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08321__C _01658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10423__I _04308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10061_ _04148_ mod.u_cpu.rf_ram.memory\[508\]\[0\] _04152_ _04153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_134_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_251_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_229_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13820_ _06311_ _06458_ _06466_ _06372_ _06776_ _06819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_169_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_251_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07732__I _01444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13751_ _06323_ _06425_ _06326_ _06281_ _06330_ _06756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_10963_ _04719_ _04772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11520__I0 _05147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_216_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_56_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12702_ _03728_ _04643_ _05959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_141_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13682_ _06692_ _01293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_43_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10894_ _04695_ mod.u_cpu.rf_ram.memory\[378\]\[0\] _04725_ _04726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_70_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_15421_ _01196_ net3 mod.u_cpu.cpu.genblk1.align.ctrl_misal vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_54_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_12633_ _05913_ _01023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_231_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09659__I _03858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_180_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15352_ _01127_ net3 mod.u_cpu.cpu.ctrl.i_iscomp vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12564_ _05855_ mod.u_cpu.rf_ram.memory\[160\]\[0\] _05866_ _05867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_180_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_196_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14303_ _00157_ net3 mod.u_cpu.rf_ram.memory\[536\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_54_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11515_ _05147_ mod.u_cpu.rf_ram.memory\[281\]\[1\] _05150_ _05152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_200_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14803__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15283_ _00042_ net4 mod.u_scanchain_local.module_data_in\[40\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_184_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12495_ _05822_ mod.u_cpu.rf_ram.memory\[170\]\[1\] _05820_ _05823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_141_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_138_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14234_ _00088_ net3 mod.u_cpu.rf_ram.memory\[570\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11446_ _05102_ _00647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13725__B2 _06314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14165_ _03670_ _07072_ _07074_ _07075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_11377_ _05057_ _00623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_166_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_256_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13116_ _06230_ mod.u_cpu.rf_ram.memory\[0\]\[0\] _06245_ _06246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_153_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14953__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10328_ _04251_ _03886_ _04342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_14096_ _07021_ mod.u_cpu.rf_ram.memory\[120\]\[0\] _07030_ _07031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09157__A1 mod.u_arbiter.i_wb_cpu_rdt\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14150__A1 _07026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13047_ _04067_ _05387_ _06201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10259_ _04293_ _00269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_79_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_266_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_266_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07263__S0 _01567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15309__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_239_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13644__I _06655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14998_ _00852_ net3 mod.u_cpu.rf_ram.memory\[66\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_207_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12464__A1 _05790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_241_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13949_ _03438_ _06917_ _06919_ _06922_ _06923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_235_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_235_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08132__A2 _02439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14333__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_207_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07470_ _01757_ _01778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_35_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__15459__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15619_ _01390_ net3 mod.u_cpu.rf_ram.memory\[247\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_195_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09140_ _03433_ _03434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_203_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09632__A2 _03837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_198_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__14483__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07643__A1 _01949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09071_ _03372_ _03373_ _03374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_120_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08022_ mod.u_cpu.rf_ram.memory\[119\]\[0\] _02330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_129_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13567__I1 mod.u_arbiter.i_wb_cpu_dbus_adr\[18\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_200_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_190_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_235_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07817__I _01672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09973_ _04091_ mod.u_cpu.rf_ram.memory\[522\]\[1\] _04088_ _04092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_131_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11339__I _05031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5009 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08924_ _02534_ _03230_ _03231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_170_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09943__I0 _04071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08855_ _03017_ _03154_ _03161_ _02852_ _03162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_258_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_218_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08371__A2 _02667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07806_ _02111_ mod.u_cpu.rf_ram.memory\[172\]\[0\] _02113_ _02114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_3629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08786_ mod.u_cpu.rf_ram.memory\[88\]\[1\] mod.u_cpu.rf_ram.memory\[89\]\[1\] mod.u_cpu.rf_ram.memory\[90\]\[1\]
+ mod.u_cpu.rf_ram.memory\[91\]\[1\] _01673_ _01855_ _03093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_73_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_233_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2906 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_226_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2917 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2928 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07737_ _02040_ _02044_ _02045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_2939 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_214_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_198_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07668_ _01739_ _01944_ _01975_ _01976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_25_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_214_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09407_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[28\] _03642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_111_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14826__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_201_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07599_ _01663_ _01906_ _01907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_200_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15421__D _01196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10069__I0 _04157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_213_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_205_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09338_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[17\] _03583_ _03584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_16_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_178_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07634__A1 _01918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09269_ _03524_ _03525_ _03526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_11300_ _05005_ _00598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__14976__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13558__I1 mod.u_arbiter.i_wb_cpu_dbus_adr\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12280_ _05428_ _05668_ _05672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11231_ mod.u_cpu.rf_ram.memory\[325\]\[0\] _04954_ _04956_ _04957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__13183__A2 mod.u_arbiter.i_wb_cpu_rdt\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_84_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11162_ _04766_ _04906_ _04910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_121_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07493__S0 _01753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11249__I _04905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10792__I1 mod.u_cpu.rf_ram.memory\[394\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14132__A1 _03850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10113_ _03842_ _04189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_136_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11093_ _04863_ _00533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_5521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_49_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_49_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_212_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09934__I0 _04054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10044_ _04140_ mod.u_cpu.rf_ram.memory\[511\]\[1\] _04138_ _04141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_14921_ _00775_ net3 mod.u_cpu.rf_ram.memory\[149\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_5554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_102_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_5587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_248_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14356__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14852_ _00706_ net3 mod.u_cpu.rf_ram.memory\[261\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_91_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07462__I _01741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15601__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_264_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4897 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13803_ _06424_ _06803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_95_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_223_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14783_ _00637_ net3 mod.u_cpu.rf_ram.memory\[296\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_21_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11995_ _05464_ mod.u_cpu.rf_ram.memory\[569\]\[1\] _05478_ _05480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_16_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_217_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_232_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13734_ _06723_ mod.u_arbiter.i_wb_cpu_rdt\[17\] _06740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__12997__A2 _03404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_189_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_188_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10946_ _04761_ _00488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_232_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14199__A1 _03389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13665_ _06338_ _06659_ _06665_ _06676_ _06677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_71_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_220_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10877_ _04611_ _04714_ _04715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__11712__I _05254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_262_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12749__A2 _05989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15404_ _01179_ net3 mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_31_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_12616_ _05902_ _01017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13596_ mod.u_arbiter.i_wb_cpu_dbus_adr\[30\] _03694_ _06619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_197_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__09614__A2 _03823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15335_ _01110_ net3 mod.u_cpu.rf_ram.memory\[89\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_200_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12547_ _05649_ _05831_ _05856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11421__A2 _05085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15266_ _00023_ net4 mod.u_arbiter.i_wb_cpu_rdt\[21\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_172_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12478_ _05811_ _00970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_172_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14217_ _04025_ _05263_ _07106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11429_ _05087_ mod.u_cpu.rf_ram.memory\[294\]\[1\] _05090_ _05092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_160_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10264__S _04295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15197_ _01050_ net3 mod.u_cpu.rf_ram.memory\[7\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_153_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07928__A2 mod.u_cpu.rf_ram.memory\[228\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10232__I0 _04267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08050__A1 _01823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14148_ _07063_ _01388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07484__S0 _01745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09057__C _03359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_258_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15131__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14079_ _07019_ _01363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_100_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input5_I io_in[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08896__C _02489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_79_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09550__A1 _03767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08640_ _02130_ _02946_ _02947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_66_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_227_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15281__CLK net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07372__I _01679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_215_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08571_ _01962_ mod.u_cpu.rf_ram.memory\[276\]\[1\] _02877_ _02878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_82_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12437__A1 _05325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14849__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08105__A2 _02412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_07522_ _01820_ _01830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_81_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08656__A3 _02962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_179_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_223_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07453_ _01759_ _01760_ _01761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11622__I _05221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14999__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_195_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07384_ _01678_ _01685_ _01691_ _01692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_206_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11799__I0 _05342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09123_ _03362_ _03385_ _03421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_191_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_176_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09054_ _03356_ _03357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_194_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_191_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__14229__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08005_ mod.u_cpu.rf_ram.memory\[125\]\[0\] _02313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__09369__A1 _03568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08416__I0 mod.u_cpu.rf_ram.memory\[408\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_191_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12212__I1 _05617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_237_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07919__A2 mod.u_cpu.rf_ram.memory\[212\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_144_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10923__A1 _04184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09956_ _04080_ _00179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__14379__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__15624__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08907_ _02525_ _03210_ _03213_ _02467_ _03214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_4105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_106_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_264_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09887_ _03995_ _04033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_4127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08838_ mod.u_cpu.rf_ram.memory\[56\]\[1\] mod.u_cpu.rf_ram.memory\[57\]\[1\] mod.u_cpu.rf_ram.memory\[58\]\[1\]
+ mod.u_cpu.rf_ram.memory\[59\]\[1\] _02242_ _02388_ _03145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_3404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_218_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12428__A1 _05759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_205_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08769_ _02283_ _03072_ _03075_ _02308_ _03076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_260_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_199_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10800_ _04531_ _04661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_2747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_226_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_214_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11780_ _05311_ mod.u_cpu.rf_ram.memory\[235\]\[0\] _05331_ _05332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_2769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10731_ _04598_ mod.u_cpu.rf_ram.memory\[404\]\[0\] _04614_ _04615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_81_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07855__A1 _01819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_214_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_207_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_186_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_202_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15004__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_201_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_13450_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[9\] _06525_ _06526_ _03541_ _06528_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_90_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10662_ _03993_ _04132_ _04568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_201_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09002__I _01430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12401_ _05695_ _05753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_51_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_222_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11403__A2 _05058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13381_ _06413_ _06461_ _06474_ _06476_ _06477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_16_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12564__S _05866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10593_ _04521_ _00375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_194_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15120_ _00973_ net3 mod.u_cpu.rf_ram.memory\[171\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12332_ _05706_ _00929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_194_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_166_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__15154__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15051_ _00905_ net3 mod.u_cpu.rf_ram.memory\[194\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12263_ _05634_ _05660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_181_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14002_ _06963_ _06964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07457__I _01527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11214_ _04944_ _00573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_123_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12194_ _05613_ _00884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_162_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14105__A1 _03836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11145_ mod.u_cpu.rf_ram.memory\[33\]\[0\] _04658_ _04898_ _04899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_150_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_5340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11076_ _03750_ _04852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_49_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11714__I0 _05268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10517__I1 mod.u_cpu.rf_ram.memory\[440\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09532__A1 _03753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08335__A2 _02637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14904_ _00758_ net3 mod.u_cpu.rf_ram.memory\[232\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_209_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10027_ mod.u_cpu.rf_ram.memory\[513\]\[1\] _04111_ _04126_ _04128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_5384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_209_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07192__I _01499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10142__A2 _04202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_263_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11190__I1 mod.u_cpu.rf_ram.memory\[332\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_252_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14835_ _00689_ net3 mod.u_cpu.rf_ram.memory\[270\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_224_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_184_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3960 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11643__S _05236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3971 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3982 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3993 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14766_ _00620_ net3 mod.u_cpu.rf_ram.memory\[304\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_189_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11978_ mod.u_cpu.rf_ram.memory\[549\]\[1\] _05468_ _05466_ _05469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_45_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_229_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09835__A2 _03996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_220_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13717_ _06723_ mod.u_arbiter.i_wb_cpu_rdt\[16\] _06724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10929_ _03841_ _04749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__11642__A2 _04026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14697_ _00551_ net3 mod.u_cpu.rf_ram.memory\[33\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_108_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13919__A1 _03403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13648_ _06289_ _06313_ _06361_ _06393_ _06660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_158_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_220_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_192_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13395__A2 _06329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13579_ mod.u_arbiter.i_wb_cpu_dbus_adr\[22\] mod.u_arbiter.i_wb_cpu_dbus_adr\[23\]
+ _06609_ _06610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_201_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_200_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08271__A1 _02550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15318_ _01097_ net3 mod.u_cpu.raddr\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_117_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_68_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__13369__I _06464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_195_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12273__I _05666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_195_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15249_ _00074_ net4 mod.u_arbiter.i_wb_cpu_rdt\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_114_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_236_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14521__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10205__I0 _04249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08023__A1 _01863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10756__I1 mod.u_cpu.rf_ram.memory\[400\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_259_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09810_ _03977_ _00136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_154_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08574__A2 mod.u_cpu.rf_ram.memory\[278\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_45_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09741_ _03696_ _03923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_246_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__14671__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09523__A1 _03271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09672_ _03862_ mod.u_cpu.rf_ram.memory\[561\]\[1\] _03867_ _03869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09523__B2 _01461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_228_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08623_ mod.u_cpu.rf_ram.memory\[156\]\[1\] mod.u_cpu.rf_ram.memory\[157\]\[1\] mod.u_cpu.rf_ram.memory\[158\]\[1\]
+ mod.u_cpu.rf_ram.memory\[159\]\[1\] _01925_ _02071_ _02930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_215_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_242_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15027__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08554_ _01938_ mod.u_cpu.rf_ram.memory\[318\]\[1\] _02860_ _01952_ _02861_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__12130__I0 _05559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07505_ _01770_ _01801_ _01811_ _01812_ _01813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_223_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07837__A1 _02105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_211_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08485_ mod.u_cpu.rf_ram.memory\[359\]\[1\] _02792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_126_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12830__A1 _03781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07436_ _01743_ _01744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_126_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_211_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_202_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15177__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13386__A2 _06447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07367_ _01670_ _01674_ _01675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_148_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_182_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09757__I _03889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09106_ _03398_ mod.u_cpu.cpu.state.ibus_cyc _03406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_182_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07298_ mod.u_cpu.rf_ram.memory\[504\]\[0\] mod.u_cpu.rf_ram.memory\[505\]\[0\] mod.u_cpu.rf_ram.memory\[506\]\[0\]
+ mod.u_cpu.rf_ram.memory\[507\]\[0\] _01605_ _01570_ _01606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_191_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_191_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13279__I _06116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12183__I _05604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09037_ _03337_ _03339_ _03340_ _03341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_201_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_163_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_85_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08014__A1 _02293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08565__A2 _02864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09762__A1 _03818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_266_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_266_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_213_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09939_ _04033_ _04068_ _04069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_265_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12950_ _06116_ mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat\[1\] _06127_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13310__A2 _06407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_219_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_133_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_219_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_245_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_234_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11901_ _05406_ mod.u_cpu.rf_ram.memory\[225\]\[1\] _05414_ _05416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_3223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12881_ _03968_ _06048_ _06077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_206_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_22_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_234_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_261_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11832_ _05310_ _05366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_3278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14620_ _00474_ net3 mod.u_cpu.rf_ram.memory\[377\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_199_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_214_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14551_ _00405_ net3 mod.u_cpu.rf_ram.memory\[412\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11763_ _05252_ _05319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_1854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10714_ _04542_ _04603_ _04604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_13502_ _03648_ _06557_ _06558_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[30\] _06560_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__13898__B _06847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14482_ _00336_ net3 mod.u_cpu.rf_ram.memory\[446\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1898 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11694_ _05272_ _00725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__14023__B1 _06971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_220_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__13377__A2 _06464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13433_ _06517_ _01219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_10645_ _04522_ _04557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_167_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14544__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13364_ _06422_ _06459_ _06460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_155_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_194_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10576_ _04510_ _00369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_127_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15103_ _00957_ net3 mod.u_cpu.rf_ram.memory\[489\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10060__A1 _03782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12315_ _05694_ _05695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_255_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__14225__D _00001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10606__I _03733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_181_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13295_ _06392_ _06393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_170_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07187__I _01494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15034_ _00888_ net3 mod.u_cpu.rf_ram.memory\[200\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_154_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_218_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12246_ _05648_ _00901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_181_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_218_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_181_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14694__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08556__A2 _02855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12177_ _05325_ _05568_ _05601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_155_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_257_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11128_ _04741_ _04887_ _04888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_228_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11059_ _04838_ _04704_ _04839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_5181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_225_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_266_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11863__A2 _05388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_225_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_224_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_266_1349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__14101__I1 mod.u_cpu.rf_ram.memory\[110\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14818_ _00672_ net3 mod.u_cpu.rf_ram.memory\[278\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_149_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08746__I mod.u_cpu.rf_ram.memory\[109\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_251_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_240_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07650__I _01827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09808__A2 _03975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14749_ _00603_ net3 mod.u_cpu.rf_ram.memory\[313\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12812__A1 _04844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_178_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09284__A3 _03521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_264_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_220_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08270_ _02139_ _02578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_32_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_220_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_165_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07221_ _01528_ _01529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_193_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_203_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_192_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11379__A1 _04775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07152_ _01460_ _01461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_157_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09744__A1 _03714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12731__I _05919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11551__A1 _04758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_232_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_247_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07985_ _01669_ _02293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_101_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11347__I _03849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09724_ _03909_ _03910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_210_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_132_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_228_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_227_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_216_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_210_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09655_ _03757_ _03855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__14417__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_243_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_216_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_216_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08606_ _01470_ _02836_ _02912_ _02913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_167_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09586_ _03800_ mod.u_cpu.rf_ram.memory\[570\]\[1\] _03798_ _03801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08537_ mod.u_cpu.rf_ram.memory\[288\]\[1\] mod.u_cpu.rf_ram.memory\[289\]\[1\] mod.u_cpu.rf_ram.memory\[290\]\[1\]
+ mod.u_cpu.rf_ram.memory\[291\]\[1\] _01826_ _02164_ _02844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_208_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_196_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_243_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14567__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08483__A1 _01520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08468_ _01855_ _02771_ _02774_ _01631_ _02775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_169_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_196_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07419_ _01705_ mod.u_cpu.rf_ram.memory\[404\]\[0\] _01726_ _01727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_196_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08399_ mod.u_cpu.rf_ram.memory\[439\]\[1\] _02706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_177_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09487__I _03712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10430_ _04106_ _04412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_137_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10361_ _04347_ _04365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_191_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_192_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_191_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12100_ _05404_ _05549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_151_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13080_ _06222_ _01161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_163_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10292_ _04318_ _00277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_88_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_219_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_152_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11458__S _05111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12031_ _05504_ _00830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12641__I _05886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_239_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_266_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_144_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_77_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13982_ mod.u_arbiter.i_wb_cpu_dbus_dat\[9\] _06943_ _06949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_92_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11145__I1 _04658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3020 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_234_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3031 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12933_ _06062_ _03669_ _06111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_207_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_206_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3042 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15342__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_248_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3053 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3064 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13047__A1 _04067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3075 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_233_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_12864_ _06064_ _06065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3086 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_222_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07470__I _01757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3097 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14603_ _00457_ net3 mod.u_cpu.rf_ram.memory\[386\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_261_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11815_ _03949_ _05355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_61_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13598__A2 _03669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15583_ _01354_ net3 mod.u_arbiter.i_wb_cpu_dbus_dat\[25\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12795_ _06020_ _01078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_226_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_202_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11746_ _02412_ _05306_ _05307_ _00742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__08474__A1 _01729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__15492__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14534_ _00388_ net3 mod.u_cpu.rf_ram.memory\[420\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_187_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_230_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_186_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_175_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11677_ _05260_ _00720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_169_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14465_ _00319_ net3 mod.u_cpu.rf_ram.memory\[455\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_70_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08515__B _02821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_174_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10628_ _04537_ mod.u_cpu.rf_ram.memory\[422\]\[1\] _04545_ _04547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_13416_ _06505_ _01214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_14396_ _00250_ net3 mod.u_cpu.rf_ram.memory\[48\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_259_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13347_ _06442_ _06314_ _06443_ _06382_ _06444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_143_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10336__I _04347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_183_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10559_ _04499_ _00363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_142_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10584__A2 _04507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_182_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13278_ _06306_ _06364_ _06370_ _06372_ _06375_ _06376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_154_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09726__A1 _03902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15017_ _00871_ net3 mod.u_cpu.rf_ram.memory\[207\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12229_ _05226_ _05594_ _05637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_142_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_96_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08250__B _01447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_190_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_233_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_233_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_229_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11167__I _04067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_256_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07770_ _02065_ _02069_ _02073_ _02076_ _02077_ _02078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_68_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09860__I _03836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_209_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08701__A2 _03004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09440_ _03395_ _03331_ _03671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_92_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_266_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__14086__I0 _06904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07380__I _01687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_225_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_213_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09371_ _03610_ _03608_ _03611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_80_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10647__I0 _04557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08322_ _02609_ _02619_ _02628_ _02629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_221_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07268__A2 mod.u_cpu.rf_ram.memory\[468\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_240_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10272__A1 _04299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08253_ _02107_ _02561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_166_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_193_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09009__A3 _03260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07204_ mod.u_cpu.rf_ram.memory\[453\]\[0\] _01512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__13210__A1 _06309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08184_ _02471_ _02474_ _02490_ _02491_ _02492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_118_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10024__A1 _04125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11072__I0 _04843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07135_ _01419_ _01443_ _01444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_161_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_238_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11772__A1 _05325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15215__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10182__S _04239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_245_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08076__S0 _02366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07555__I _01862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_1246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15365__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_199_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_114_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08587__S _02106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07968_ _02174_ _02271_ _02275_ _01766_ _02276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__13277__A1 _06321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09707_ _03893_ _03896_ _03897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__11827__A2 _05362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07899_ _01787_ _02207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_67_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_74_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_249_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09638_ _03841_ _03842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_215_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_167_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_204_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08319__C _01751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09569_ _03700_ _03743_ _03787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_43_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_231_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_231_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11600_ _05207_ _00696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_208_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_169_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10638__I0 _04537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12580_ _05874_ mod.u_cpu.rf_ram.memory\[158\]\[1\] _05876_ _05878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08456__A1 _02711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_180_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_211_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_208_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11531_ _05107_ _05162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_212_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10263__A1 _02439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14250_ _00104_ net3 mod.u_cpu.rf_ram.memory\[562\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_184_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11462_ _05045_ _05114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_184_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12004__A2 _04984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_137_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_11_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09010__I _01428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13201_ _06302_ _06303_ _06308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__08054__C _02361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11063__I0 _04841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10413_ _04255_ _04373_ _04401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_109_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14181_ _07085_ _01399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08303__S1 _02454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_256_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_11393_ _05068_ _00628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_165_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09945__I _04050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13132_ mod.u_arbiter.i_wb_cpu_rdt\[18\] mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat\[2\]
+ _06253_ _06256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_178_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10344_ _04352_ _04353_ _04354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_87_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13467__I _06537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_174_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13063_ _06211_ _01155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10275_ _04288_ mod.u_cpu.rf_ram.memory\[478\]\[1\] _04304_ _04306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_191_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10318__A2 _04335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07465__I _01750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12014_ _05484_ mod.u_cpu.rf_ram.memory\[57\]\[1\] _05491_ _05493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_65_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_215_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_238_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13268__A1 _06318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14732__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_266_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13965_ mod.u_arbiter.i_wb_cpu_dbus_dat\[5\] _06917_ _06918_ _06935_ _06936_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_171_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_262_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12916_ mod.u_cpu.rf_ram.memory\[389\]\[0\] _05971_ _06099_ _06100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_73_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13896_ _06884_ _01315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_46_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12491__A2 _05767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15635_ _01406_ net3 mod.u_cpu.cpu.state.o_cnt_r\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__14882__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_222_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12847_ _02080_ _03742_ _06053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_2171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_261_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_250_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11651__S _05240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_222_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_203_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08447__A1 _02230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15566_ _01337_ net3 mod.u_arbiter.i_wb_cpu_dbus_dat\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12778_ _06008_ _01073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_159_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_222_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_187_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14517_ _00371_ net3 mod.u_cpu.rf_ram.memory\[42\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11729_ _05287_ mod.u_cpu.rf_ram.memory\[242\]\[1\] _05294_ _05296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_147_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13991__A2 _06952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_175_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11450__I _03732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15497_ _01268_ net3 mod.u_arbiter.i_wb_cpu_dbus_adr\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_187_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15238__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_174_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14448_ _00302_ net3 mod.u_cpu.rf_ram.memory\[463\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_80_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_200_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_174_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13743__A2 _06456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14379_ _00233_ net3 mod.u_cpu.rf_ram.memory\[498\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_183_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14262__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15388__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11098__S _04865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08940_ _01466_ _02914_ _03167_ _03246_ _00001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_170_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12554__I0 _05855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08871_ mod.u_cpu.rf_ram.memory\[557\]\[1\] _03178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_97_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07308__C _01615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07822_ _01744_ _02130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08922__A2 mod.u_cpu.rf_ram.memory\[540\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_257_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13259__A1 _05787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09590__I _03803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12306__I0 _05677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_226_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07753_ _02057_ _02060_ _01632_ _02061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_226_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14001__I _05801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07684_ _01991_ _01992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_38_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07489__A2 _01796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_252_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_198_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09423_ _03564_ _03655_ _03656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_53_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_213_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_244_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_240_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09354_ _03597_ _00060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__12234__A2 _04227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_178_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08305_ mod.u_cpu.rf_ram.memory\[477\]\[1\] _02612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_21_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09285_ mod.u_cpu.cpu.ctrl.o_ibus_adr\[9\] _03538_ _03539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__07110__A1 _01418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11360__I _05045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_166_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08236_ mod.u_cpu.rf_ram.memory\[520\]\[0\] mod.u_cpu.rf_ram.memory\[521\]\[0\] mod.u_cpu.rf_ram.memory\[522\]\[0\]
+ mod.u_cpu.rf_ram.memory\[523\]\[0\] _02507_ _02543_ _02544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_53_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11045__I0 _04825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14605__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_193_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13734__A2 mod.u_arbiter.i_wb_cpu_rdt\[17\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08167_ _01702_ _02475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_107_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07118_ mod.u_cpu.cpu.decode.op21 _01426_ _01427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_88_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08098_ _01644_ _02406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__07413__A2 _01699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08602__C _01887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12191__I _05432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14755__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10060_ _03782_ _04143_ _04152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_216_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07218__C _01525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_248_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09206__S _03474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_217_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_244_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13750_ _03510_ mod.u_arbiter.i_wb_cpu_rdt\[18\] _06754_ _06755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08677__A1 _02462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10962_ _01897_ _04770_ _04771_ _00494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_84_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__13670__A1 _06651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_189_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12701_ _05958_ _01046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_252_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_243_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13681_ mod.u_cpu.cpu.immdec.imm19_12_20\[1\] _06691_ _06658_ _06692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_10893_ _04322_ _04709_ _04725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_232_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15420_ _01195_ net3 mod.u_cpu.rf_ram.memory\[349\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_12632_ _05904_ mod.u_cpu.rf_ram.memory\[14\]\[0\] _05912_ _05913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_19_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08429__A1 _02534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__13422__A1 _03377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_262_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10236__A1 _04277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15351_ _01126_ net3 mod.u_cpu.cpu.genblk3.csr.o_new_irq vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12563_ _05417_ _05757_ _05866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__11270__I _04844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_157_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11514_ _05151_ _00666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_157_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14302_ _00156_ net3 mod.u_cpu.rf_ram.memory\[536\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_7_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12494_ _05806_ _05822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_15282_ _00040_ net4 mod.u_scanchain_local.module_data_in\[39\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__14285__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_221_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11036__I0 _04803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14233_ _00087_ net3 mod.u_cpu.rf_ram.memory\[571\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11445_ _05087_ mod.u_cpu.rf_ram.memory\[291\]\[1\] _05100_ _05102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_144_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15530__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08288__S0 _02593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12784__I0 _06010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14164_ _03298_ _07073_ _07074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_11376_ _05050_ mod.u_cpu.rf_ram.memory\[303\]\[1\] _05055_ _05057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08601__A1 _02323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13115_ _06181_ _03986_ _06245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_152_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10327_ _04341_ _00289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_152_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14095_ _03804_ _07014_ _07030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_152_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09157__A2 _03436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13046_ _06200_ _01149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_10258_ _04288_ mod.u_cpu.rf_ram.memory\[480\]\[1\] _04291_ _04293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_59_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07168__A1 _01447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_239_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_227_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07263__S1 _01570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10189_ _04244_ _00248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_113_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14997_ _00851_ net3 mod.u_cpu.rf_ram.memory\[65\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_47_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_208_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08668__A1 _01567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13948_ _06920_ _06921_ _06922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__13661__A1 _06309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_234_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_207_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_263_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_13879_ mod.u_arbiter.i_wb_cpu_rdt\[24\] mod.u_arbiter.i_wb_cpu_rdt\[8\] _06334_
+ _06871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_61_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_222_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15618_ _01389_ net3 mod.u_cpu.rf_ram.memory\[247\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__15060__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_98_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_203_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14628__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15549_ _01320_ net3 mod.u_cpu.cpu.decode.co_mem_word vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_72_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11975__A1 _05322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09070_ _01434_ _01436_ _03373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__14213__I0 _03699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_175_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08021_ _02134_ _02329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_163_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_200_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14778__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08703__B _01891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_190_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_239_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08422__C _01773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12940__S _06116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09972_ _04090_ _04091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_143_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08923_ mod.u_cpu.rf_ram.memory\[543\]\[1\] _03230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_131_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07159__A1 _01463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_130_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08854_ _02063_ _03157_ _03160_ _01695_ _03161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_131_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07805_ _01673_ _02112_ _02113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_3619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08785_ _01696_ _03091_ _01720_ _03092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_85_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_211_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2907 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07736_ mod.u_cpu.rf_ram.memory\[128\]\[0\] mod.u_cpu.rf_ram.memory\[129\]\[0\] mod.u_cpu.rf_ram.memory\[130\]\[0\]
+ mod.u_cpu.rf_ram.memory\[131\]\[0\] _02041_ _02043_ _02044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_2918 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15403__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2929 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_253_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_198_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07667_ _01740_ _01955_ _01974_ _01975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_246_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_225_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_214_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11291__S _04997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09406_ _03623_ _03640_ _03641_ _00069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_198_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_40_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_241_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13404__A1 _06483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07598_ mod.u_cpu.rf_ram.memory\[359\]\[0\] _01906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_213_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11266__I0 _04976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_90_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_231_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_166_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15553__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09337_ _03582_ _03579_ _03583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_194_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09268_ _03520_ _03521_ _03525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__08831__A1 _02405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_194_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11018__I0 _04797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08219_ _02526_ _02527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13707__A2 _06667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09199_ mod.u_arbiter.i_wb_cpu_rdt\[25\] mod.u_arbiter.i_wb_cpu_dbus_dat\[22\] _03469_
+ _03472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_147_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12766__I0 _05992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11230_ _04955_ _04922_ _04956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_140_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12391__A1 _03770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11161_ _04909_ _00555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_122_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07493__S1 _01771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12518__I0 _05837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10112_ _04188_ _00227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_150_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__14132__A2 _05631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11092_ _04862_ mod.u_cpu.rf_ram.memory\[348\]\[1\] _04860_ _04863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_249_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_216_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_251_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10043_ _04090_ _04140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_14920_ _00774_ net3 mod.u_cpu.rf_ram.memory\[149\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_121_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09444__B _03674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08442__S0 _02020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_212_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07743__I _01661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14851_ _00705_ net3 mod.u_cpu.rf_ram.memory\[262\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_5599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07570__A1 _01875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_236_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13802_ _06418_ _06466_ _06666_ _06443_ _06486_ _06802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_5_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__15083__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4898 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_205_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_14782_ _00636_ net3 mod.u_cpu.rf_ram.memory\[296\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__13643__A1 _03390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_217_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11994_ _05479_ _00818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_216_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13733_ _06723_ _06739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_10945_ _04753_ mod.u_cpu.rf_ram.memory\[370\]\[0\] _04760_ _04761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_205_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13664_ _06672_ _06674_ _06675_ _06472_ _06134_ _06676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_10876_ _04307_ _04713_ _04714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__10209__A1 _03942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_227_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_220_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11257__I0 _04961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15403_ _01178_ net3 mod.u_cpu.cpu.genblk1.align.ibus_rdt_concat\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08507__C _02453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_231_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_188_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_12615_ _05887_ mod.u_cpu.rf_ram.memory\[152\]\[0\] _05901_ _05902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XPHY_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_13595_ _06618_ _01280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_185_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15334_ _01109_ net3 mod.u_cpu.rf_ram.memory\[99\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08822__A1 _02405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14920__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12546_ _05812_ _05855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_200_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15265_ _00022_ net4 mod.u_arbiter.i_wb_cpu_rdt\[20\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12477_ _05807_ mod.u_cpu.rf_ram.memory\[519\]\[1\] _05809_ _05811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_8_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12757__I0 _05984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14216_ _07105_ _01415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_67_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11428_ _05091_ _00640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_15196_ _01049_ net3 mod.u_cpu.rf_ram.memory\[7\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_99_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_158_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10232__I1 mod.u_cpu.rf_ram.memory\[484\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11359_ _04959_ _05045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_153_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12760__S _05996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14147_ _07055_ mod.u_cpu.rf_ram.memory\[90\]\[1\] _07061_ _07063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_152_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_193_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07484__S1 _01747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_180_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14078_ _06578_ mod.u_cpu.rf_ram.memory\[299\]\[0\] _07018_ _07019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12134__A1 _05334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11376__S _05055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13029_ _06189_ _01143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_112_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__14300__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13882__A1 _06858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15426__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09550__A2 _03771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_120_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07561__A1 _01855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08570_ _01963_ _02876_ _02877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_148_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12437__A2 _05767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_254_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_235_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07521_ mod.u_cpu.rf_ram.memory\[328\]\[0\] mod.u_cpu.rf_ram.memory\[329\]\[0\] mod.u_cpu.rf_ram.memory\[330\]\[0\]
+ mod.u_cpu.rf_ram.memory\[331\]\[0\] _01826_ _01828_ _01829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__10448__A1 _04281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_223_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_207_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15576__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14450__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11903__I _03984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07452_ mod.u_cpu.rf_ram.memory\[423\]\[0\] _01760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_22_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_228_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07321__C _01587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07383_ _01688_ _01690_ _01691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_188_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09122_ _03363_ _03416_ _03420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_163_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_241_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_198_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09053_ _03308_ _03356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_159_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07828__I _01862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08004_ mod.u_cpu.rf_ram.memory\[120\]\[0\] mod.u_cpu.rf_ram.memory\[121\]\[0\] mod.u_cpu.rf_ram.memory\[122\]\[0\]
+ mod.u_cpu.rf_ram.memory\[123\]\[0\] _02294_ _02295_ _02312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_159_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10254__I _03985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10923__A2 _04713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09955_ mod.u_cpu.rf_ram.memory\[525\]\[1\] _03929_ _04078_ _04080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_106_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13322__B1 _06339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08906_ _02533_ mod.u_cpu.rf_ram.memory\[518\]\[1\] _03212_ _02537_ _03213_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_253_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13873__A1 _06739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09886_ _04032_ _00157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_258_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_170_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_106_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_218_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_4128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_170_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08837_ mod.u_cpu.rf_ram.memory\[60\]\[1\] mod.u_cpu.rf_ram.memory\[61\]\[1\] mod.u_cpu.rf_ram.memory\[62\]\[1\]
+ mod.u_cpu.rf_ram.memory\[63\]\[1\] _02406_ _02218_ _03144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_3405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07552__A1 _01858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08768_ _02316_ mod.u_cpu.rf_ram.memory\[126\]\[1\] _03074_ _02306_ _03075_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_2715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07719_ _02026_ _02027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_54_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13514__B _03337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12979__A3 _06153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_214_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_199_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08699_ _02190_ _03005_ _03006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_25_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_214_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_198_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_198_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10730_ _04189_ _04599_ _04614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__07855__A2 _02162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__14943__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_213_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11239__I0 _04961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09057__A1 _03355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10661_ _04567_ _00397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_186_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_41_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12400_ _05752_ _00951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_210_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13380_ _06139_ _06475_ _06476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08804__A1 _01511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10592_ _04514_ mod.u_cpu.rf_ram.memory\[427\]\[1\] _04519_ _04521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09852__I0 _03999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_194_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10611__A1 _04255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12331_ _05692_ mod.u_cpu.rf_ram.memory\[184\]\[1\] _05704_ _05706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_215_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_177_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12262_ _05659_ _00906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_15050_ _00904_ net3 mod.u_cpu.rf_ram.memory\[194\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_108_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09604__I0 _03802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_182_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11213_ _04936_ mod.u_cpu.rf_ram.memory\[328\]\[1\] _04942_ _04944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_141_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14001_ _05801_ _06963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_257_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput6 net6 io_out[13] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_181_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12193_ _05605_ mod.u_cpu.rf_ram.memory\[202\]\[0\] _05612_ _05613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__14323__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__15449__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11144_ _03809_ _03980_ _04898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__14105__A2 _05720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12116__A1 _05293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13313__B1 _06400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11075_ _04851_ _00527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_163_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13864__A1 _06856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12911__I0 _06088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14903_ _00757_ net3 mod.u_cpu.rf_ram.memory\[233\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_114_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10026_ _04127_ _00202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_5374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_248_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_188_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09532__A2 _03755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__14473__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__15599__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_209_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14834_ _00688_ net3 mod.u_cpu.rf_ram.memory\[270\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_4673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_264_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13616__A1 _06249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3950 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_236_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3961 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_217_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3972 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14765_ _00619_ net3 mod.u_cpu.rf_ram.memory\[305\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_205_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3983 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3994 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11977_ _05229_ _05468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_45_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_264_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_225_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13716_ _05784_ _06723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_10928_ _04748_ _00483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_260_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14696_ _00550_ net3 mod.u_cpu.rf_ram.memory\[33\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_147_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_232_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_189_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_232_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_176_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13647_ mod.u_arbiter.i_wb_cpu_rdt\[20\] mod.u_arbiter.i_wb_cpu_rdt\[4\] _06334_
+ _06659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_31_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__12755__S _05993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09048__A1 _03250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10859_ mod.u_cpu.cpu.immdec.imm11_7\[3\] _04222_ _03724_ _04701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_158_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_158_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_13578_ _03692_ _06609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_121_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10602__A1 _03892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15317_ _01096_ net3 mod.u_cpu.rf_ram_if.rtrig0 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12529_ _05837_ mod.u_cpu.rf_ram.memory\[469\]\[1\] _05842_ _05845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_157_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07648__I _01914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15248_ _00063_ net4 mod.u_arbiter.i_wb_cpu_rdt\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_160_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08023__A2 _02330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15179_ _01032_ net3 mod.u_cpu.rf_ram.memory\[145\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09220__A1 _03410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_193_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_207_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14816__CLK net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13155__I0 mod.u_arbiter.i_wb_cpu_rdt\[28\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08700__C _02212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09740_ _03922_ _00121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_100_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
.ends

